PK   VH�X`C���  D�     cirkitFile.json�][��8��+��Y���T��e6��Np���DM��c���$�A��!�Kےh���Nv��`b��b��X�*�O�ƾw��rٸ���Y͖����ɽm���)�Nf�������>�On>��������w˅[��Hie��ʂ�L�Fd��6����Dߑ�͛��g�S9ÑsO>DljŤ�e&
F2�T�咹,YW�z�v�r��ͨ�rϠ6Y��(��UL;^Y?j��E�5qJeEe|�����\�9a�;^s�b��𜕪Ȍ.����(��ܕ���2�b2s�l�3�$�e�3S���Xe/�(|�����f��e�e�x���p��8r�#ϑ������شW++���X�LXM= ��\]z:n���G+��V5��:�-3P��tl����y�qYՙ0�o��E�U�%��e���i�i:�N!#&Qb#85���Bu�YR�0�Ɂ�9G�$�D�#�5��=Cnl,��H�A����H�r����.GB�ǡ[3YpAXV��[ݹ�F3��7#�������W4i!��4+%�2A5ϊ�O�ץ��V5��-
�2Ũ�ؾ��#{#�?B��s�4��K_1���u���S���5+���3 qd�ab#Z����e�Wd�1��0Tey%�m��Ǟ4�E���Z�,2Y�	iuf�1YU2!�sy�M�Ϡ�c}�|lC�d�ϕ����)
߼��<kN2MK��+�h��� �m�n$v�Ϡ�A���Ch�X����0��!�3P �gl���`�e�nmA�s���.�0`$�K�|����iԅ�E0M�a��]�C@�#��4}|c���Q�������:�C��@-ǝ+�g��h�#�Fa�����b�����4�3㞗����#R�~ޟ}����A�}N�#�߰���&�p�.�i��"6\tUD�Z���仒�G ��$㢓p1I��iP��i�K��5u^bش��k��
æ��m%0ˀ��
*<C��V*�M����P3��,�Y"�F	3���H�F�a�F�4(fiT1kQ��x��uӠ��A1OdJ�A1O�b~����w�$�[����R9�YYГ�Ӷ���s�~�t�G��\ZYr�̀H��'!^'Jq⡧g�xB�H�<Gp��P=9=r�0z�GЈ�i�B��{���F4j~u��i��>=���t.��$`���	���ǡa��04"{zt���Ӟ64RzZ�A#�	F��>F��ˠq���$4Dxڙ�F�N;�����u���W�S8m��k��-�㺱sd8υ%�pI��$\T.:	��K�u����4|i��4 �iL�@���0Mb��,�Y"��,�Y�4(fiP�Ҡ��A1K�b��<�y"S"�y�(���\��8���rVp8��,�p���9����\���Ṝ�N�s9+8���rVp8��,�p���=	N�s9+8���F��[58���rv���N� h8�����ix.gGN�s94�?O�Ǐ�Mn�ݬ�8��z:�0k���anKW��w˦r�����<y;�\N�l.����
����Z1�F�e���1�"-�,�ci������Άqc"-c^c ���d���zh|�s5cf`Z�ema������Rc,����"-��i����.�2�U���(��t$s��$����j:p��P7�0~�۷;g�q��7`Րc���ż���� /�$��%|�����pR���N
��I^8)�K�'x�/ֹ��P� /�j��z���t<�C��?.& �9)�Kx#�Sr1�����!�EI �SI �aI �oI �}�K��b�c��q��'�/��凐U�8��9�w�lb=C҇�.r�G1{��#���w��,Opr1f�4�� �s,��h�µM��hD��3�;�0} ����L"�,<���/r#�e��P�0�S��8�b��U2V'�	�(�@b`U-��a�m�,�Av�:�g��j,09�X��c��O ��џ����a�8G�9�/�H}90k8!��pA����N(�,4���.bW�S�a0�w�E�2p�1�����N"@�!�:�G�����18C�#�]_��T�s��;�ABӖ;c3����v�@7��g4������l���8w�E�/8�9�T��B��Ν��>���n ΀�Ä$\jL|q���,RprtoU}�N��̪'��W!P1S�+D���)h���0�aR�<y��i�p��Z��M;������~����
��,P�@�,P�@�Ry������
(x�Rs���ԥ�����yD �� &ڱH �� b�@l�#�vD ف� ��d�:"�h�8�C� kpǠ�T��t7�o��a��m^"�Q �d��T�[�_V�]^�ێ��m��g�٨��]q�{$�w��z�;o�_��]��Z�_l�"��vA��m|��۾��zk?� w���~�w)�o��^��q�p��}���� ���0a�%�~D�и[}�
���t�����
\�+���.�����~��!�dY��}�-ܼ�o;�=��[_�vJ趈��ض��������ĶH��H��ԶH����H��̶���mQ�+��Ѡ�����ݍ���ݍ�	�	�	ݍ�������wE�lU,mnq�˻�l�޸R�=�V?�up$?��^7�׬g����{X�
}��u3[��Z�w�{(�N���c��}+]��q1�L������/�=��Mm�+�W��m��s�ָ>�WMn�ͣ�zg��-׏�kN	pX�@�M*XI��)���z�����S}-�)��ky��l��UO��u�J)2��<S�E�d^Z[#D ����\�j���l�Z�E�e�JM'�f�؍��j�!�N9kʹ�N��ص�
J�N��y.�>�����<x����:?����<�b�SK<i-�q*�b1���|�)��Fj�y3R����:x.����#̈)g$R@",�P0�P1������X��q�78Ȝ������7�o���vP���+�Gt���UlUPR�i��W��~�m����v���[������dV�OHQ*U�U�+�Ҝ�YQ:��Fy���,�m}��a�����w�WZ�K�7�R��ʌ�$SDk"�u\�����$�Ɩ�;������m*���U�pT�J��^-��B��օΔ�,�z# ��*1Z��MW����������SO~��ͫ�N���LI�P�5ͬ�&��*��.�q�3�M�\���\��E���Rx.�.�
!|�4��TF�|�ˏ���J��Ϋ�s��8��:�s�2YV�3��:��~���]T.���mӁ[���Xl$�<���],[�Ú������Y_U�[��e��ԣON�����z�e�EX�U^R��2�
���M7-=�EU3��F�d����Y�i3�1��rB�n�S6�0a�BT<#%�2!���JI������
GX�T����D��g�ú�U&(��՚)fO#��|���_Ϊ��[?>�ן�>��.�����+�����fSrj_ݻ�M��˫�qq��{ߍ�������e4_.������ ��=8�v���Cf�usW�[̴R���d�>�������'��և�{�����]?V��~��k~�=L�6�_�����/�XU?4K[��$7����ZN3FX3�ayhOViN+�a-�QE����UT��Zy��Z���)БXמz|�YSJX�ۿ
��o�H�
?�ް}���C]�P <2�q���>v�<v2�%��l�:VU�UIP�6�f?-Z�Q�&م��� ���� �x���j�Z�0�S�v@����_R�D
�HS�������)�MO]�&��l�&��� 96���⻸��F
Vtk#�
��&h���F_4�<+ h���H;�梠�QM#.�~�r� ��l�~I���_i7�-*^��%VB��8�M^o����<���^C?��2�,�4��G4����SQmT�lF���!��D���м*E�΃�d ��u�Z4{���:,2��Bdg�G�#�"� �TC";z��d2�N��'z�Pξ�|_ٺy���^-��@�{����/E�%1�1�SNԵ��/�C��p��#�gV�i֚��pM���C���C��!^5oOL����&~��;�n_e�BJ�Ud������ ��׆I��P�A劳�ҙ_T,�����~k�N澫rx�Xg�@���4w��o�m�YI��s��\��Z*�B<K���+%��$��0��-�!F�(�k%�[��e��em�4�$*"�3��r�?2�/���#q9�lgp�]l�iz�WR�*]�*%2�ɬ�YV�FԹc��hz@�3����~���U��9T���b���#�����}A'�d���@�����j�z���$h`on���[t�G9��Idx�aV��Z9���}v��n�� �57�5M?v�8�����s��U��^����}���Nݐ��)�|ΗM{���I�����K�~=[lX�}�esL��N��]niY5�ï)E����N���l�~m��-�O�������K�:���Q����M���A�ݑYʧ���F�v�:���~��|�0:���⁐��J	
���RA�>����i���doNSN��ĉ�R  `w�@��]�b�h @��n$ ¾s�J��}G �B�����Y���v��vpH� �ҍ��.xx�J��݆���S	�'��q�%@7Ӂb��!Z*P<o� ��� ���	ƘJPk���6%(�&��ibP�00�ҍh�N���nS��!�S	�}�\CMLح_(`��[`P��n�E�N/��@%J�'|�Sk��p1b��(�;�8�%Q�t=�LӘ)W ��gy �J!���]��x����1F����uj�U�a�k�|�V{#�T��1`�{��h���9l�o$4�N��n2���]�1<�UAM�`�����؀#R�=M�:�?`-1�St`֯�uA�>�/���]�ZG^Á��; SkwTFO�]2�F!��%�'DR`�� �Ǭ�\��8�	�%�00�3j������t���?�=EeSeR�Ť�∠��R��YQ���2�3�ZhH��Zf�~1 �^�� 4B�� �s(�5z	���v+��!Z*���Hw�La�QK;�OyEcj�3��N��^����3B���G>��m����Z�ܗA�U|_
=#��z�9<��N����K�b�t_,"�BwN�@��r��޳���3B��=��k�S2S�uJ��t�'5zdRݓ=d�j�c?	T	�yL��u�Y:zL�x�l��gŉ;�a|8?5F-*��l~|�u�em+�t뢰p2��é�'�	 2��עG���!��@�� �k��*)���3�mѩ����!D�?
� kQ>�����2��EJ m��@�ퟭl� ��!�[ڋhck�&=�%����?۵kfv�����/���g�x����^�ݻ���7oV����r��[���a{sn���PK   |G�X�v��f �� /   images/153184b0-233d-45e0-a203-5756afb39f29.jpg�|w U�������JF7��\;�F$�Uff�����M������$���k�l23�M��{�T�|����߹����>��<����sn�} ͅ�
�  ���
�����������|QS�`T�h�������������	s�8�),!�/(�x����{<���e�>R"� ���}�}���� � � ���FH% ������ PB"�N F �hh  ��M.`�����l|�W�	����w���g ����v�9��Y?m$W�WV3�2�K��5�Wh�F��x����v�FI�d��UaV�k��Z��o�����
��s�g�ǆ���18��61QG6s�E̖��x�*�ގ���Rymd�2��S�zj������-S]t�8��֚:b�.�:Z���
�ޛ�]GdT��4$�I(�N�b��C�y6 �^��r�>z�W>�L;T9��u�,���&���XarEU��o��jwj��"�.y�B5�cjɩ��Cfe~�~q#�y]���e�7M9S6_Um`�\M�,_��%�ܓ��k3O��|�[�}�����K|Wf������ ��smS����~�����bw,�3{��#�I�\�m�{�SK�ĵqn���ś��j����[��Y��|�nQ�5m�q��՝�J�q�$W㞉S�<g��>.��=�A�ϣ�Ԯ��PGc�qq���bW�V��-�6=l���b#�[ b�
�;f��şx�������T����B�-k�56�#-�aK���uS�>f���w���׌�;O6�l~%�����/�Y��P��L ���k(�mx��\ �f�ጥ:F"6 Xr|�P���3���X����	�47[[*�n�J��J5�]���1�Ųo��d�wbz�#kK�Zf]��R����^z-��򴹽M{�q:hB��xe�B��t�!ͻ������n�$�[��NF����YC�����~�1f-��w���Z�+����/�5F�.*I���~~ڝ�Ʊ7��K�� S�k�c�1����Q��.$�-�@G�c�y�nx��9�Nr��D�O��D�U��x'�(���Ŷ^��B���!'-�cɝ��>��)PՅx-�
������".N��
��t�[=	O�V�?)r�!{���`�mG�`R���۰Յ=s�i��z��zw4��b�|�]�����f�0��9� ��Q��KY�7y����e%"��L�x��R��Dv�����>�۲Іy��٘"F=Qm�Qш{�L�[Ɏ�N6���KC�nW�0�/�/|��M!+iL*C[���<��g�I��ZB���Ʈ�]���ۭo��\��_ܙI:Q��T��)�;V)<r_���G#���B}2��Y9�9֚Ƶǻu���M���=�r��9��'��Kl�>�E���兄�h|��M���?�F�������J�gϟ�������/]s��D>1QS�����)��;�����G�mX��CI�o�Qˠx�?����;�����Y��G��JW���rZx'Tj�pc�H7&�`q�X�X
\�Ngy�MR�*����|��0m�	����o8FU=�6r7���5;��*����1��:w��ۀY�3��
C��#����}��K��� Z!�lЭm��"}?}r]�h9i���97��r�k��H��=�Rt\���� I�ʸ��5W��Ob�=(2d�Z�`�_���DF�8 ��PG�l�;��x��?� �}�z��x��6�^&�%�r���qA��KEk�������/��9���髃���O�6v*�
�:�?	�%�K���縹���J��[���3m f��93��{�)�zי��y���{��BW�`eR&<��B�X��3M����x�x�7�S�e_��.�w�����_��p΋B�D��۞��FJ��N�W�/:\�w?;5��N�T�|Dg�,����Q�r��b�{@��ǳ�������ht:/cafV��~>�={) �>��Dн�{�9:��|e2���B{hpF�.9�-��)x<]B<eKb���	��a{���"K�-pgڇ��';����M|(9�Uy��Q�m�8p��,��%���-�`�z��G��C{�w�)a��3w�d���h���~S�8g���F*�N=�f�"#���q��s���hD���t��N�F�>�㣌?R�N��Z6�� ���������#�>�ҷ8�uj-ݝ�sn�)�Ze�/���_v�����l#�Hi䜮wp�"�<���}kyؘhI��HU�K%h���Pp�9���(�����|�j�s.&�,�sןǲ��4K���b�t�#Z��|-�}|*$Eu-�'v4����m�y��h��:��E�k�Ln���u�y�p��Z�@P���J��z�i�3���A�[�u~��S�w��<pazsk�'>ky�j�K�ܟ%�x�x���������Bh�4�������k�o��~��f�t3��fO���c���hB���������K�?H.>_;��>I�7�hv���I�n��ec�ޒ�v����~X��C���w�y��1��Q(����8�n��P�j�pn	�[3����Y7�{q�@�D�"�{f2�Aj+�%�[Y\���Mf�V�>�m�
Ӯd.�,��8�b�=(��,.�'�$h{{m��3Ih�a9)�W%_�g�g�lk([�)��������ݴ*�h��+7;�<����9��.l�Ѡ}[t�,�e���u~ݓpș��[����y�ٳ~ұA�z��-���&�k�����	t�T�.Yn��Ng����}��O���Q쨭���W�+R9C���.���R�͢*�K����L�UY�<;��gI�#�w>[�h�E�F+=h����B�;��������[8�ώᶈc�x��&�Y�Q�ڏ!4�th.�IďǏ#� ��-<m��9�XW릢�_������=�/�|12�|�{�O|=�$�8~X45�'=�Q���vo� �4�Ϛ�l(��:�٠�C�A����Y3�H��9?	�.�<��n���P.�妗�� �}lr�R[߇ՅSw_�a���*c�1^f|���:�����X\g�wrK�����J��{ȱ��U�3&
��ܣ��\L}M�R�^�d �Փu?�ĩ+4I~{�4���F��s�����LbU$��Gn�ЅX�d�"��ʛ_s�;���N9^qmIe��f
�"�u;ʽn]��?�1� 
�=Þ�v'� ��wѡ>!�2��}w�)�Y�L��g�g�(��=+A��ؾ"TO�,22�o�Ag+��x�=]�Sh���������V*��p��u!��2^�<���pQ
�ϥ�~vY��_�T����|g�9mi��zS�Z9�wk3�}�M�/vjى�;>Rxn�Y�A�ˍ�:��`O�R��=+m���f&>ԝ�ݚ�/%��̗��`�����Оo���Vφ���wr8��;�H�ųw��-���*��qQ��"8q�����\#��pǾ�Zv����Z�2�ωt5�	�.��q������G�0��dj8Ы�{�Vd}E�:Ύ��%�~.<�赩]y�t���#�����ca'5I$��nE��+&ԒN�u>�OE���H�&_+�|w��P��Z��_py'��x>P�gP�����m^�e��Re��0����[��{\V�P.�3iA�g���7G�#O;*<;���ϭE���CK.�M����^,�3ċF�&Xr�[<6%n�ì����Lp�T{B^RN��������Ю�'�C�*?�{�W�c�<�1�[4�5z��T���T���v�w�9!�Q;E��{��$���q�� �4���!Q���y����
Z��CGl�p�n�](@��"���O�zS}Ƶ1[������mp] >�6`�b��Ȏ�y�g���^gI1���Ù�`�H�ÒK�.���j�I*�V�eJώ�9�Q�\� ���3����3�_&1q��M����� ��wz 	#w{���p����n�������ȩ|f����U�#�ΰ�����'���1zڨ5lg��M�9M���dH�"{�^�ڵ�VEvP=ͥDU��3�����u�fSݚo\��;�+�����vGQ�*.5�ՙ�5��j�m��?�H���/�v�6+N�� _M���DH�b��QE�O`�Jl�.���^��m�u��ë��++�W�������;uF3��!�G���ddZ��(wolðh������{��;8�0-g�AL�ǵ^�Uz�N���El�������#�RPv:9�2dĿ��]嵴H��b��!#h����c~���-�T��Y`�u�������-�{'������7�����2�2��DF�X���T�����t��w��"n��y6��b{��m^^ �n\s���52��#��gN>�[7δ�9��3.�M3���͛'�4�~ߓ�.�Su>(��^���x�Ģú�Y�"�l�7��W�.�AGVqt����\�qsڐ�*\�j#^*T*�3V�}ߌ�=O�V�Ix�ȵ0��;f�$[�u�GD�).ݤ�I0�k}Se�l���2�}Ҭ���4�!�^� V�ZP���f-��c�1�&1)J��$�Q���Fȥ����t���Iϲ�3x�ՏMǎ���Nގ���:8�|�F�>N�MZ��s���[SK�z��'�Jb#��1-9�/�`�;�X% ��(�$P�m�0�u�Z`^W�����'r��OO^���9�!����Y�ף�b�<�\2����������.���R����+3ײ2�����
#p�sSG�RX?��E�*��S+ �x��!h�g�����d�j�'��(� K�#W���>� ���x̽�c|;���'�z�)��r.5�"��^7��Ƭ�ާ8�Z�'2(�M��`�XN��ࠡ����n]#������\�!���:غq���
\�S��������s�*ʐ=f�Y��PJ��õZt��(�4�`K�ɍ�v�³iT͇�KÓ�<S#���K7�U�����w{�8'���/�������\��t�h��X����~�~Qͺ��ت�[H�k�'#��Z�0��*4tZ<<!q�B�ira�%���=�'cfn2u
�ȧ&(��GҏOj���k`G�]a�}�WWz�����/����y�Yh�nO�X���+r^]�q��ud{�h�^|����0Tk{�fi4��D�ِh
��bˎu�K'[�k�q�ŗF ���u�˴xt��؍���ĩ=�[]Wl;'����Ɓy�wIZoZ�҅��[m 烖n���3�H����휔���^*��1�Q1�v�lqq
�-�	Ig5��q�}P�# �k#2�m����Vy��O�.�ߩ��/��	p�8x|;6o���V՞?ݗ�n�``f���J�i�c��r,�;�]/K�7��%͎����9B��ߛ���'���-��<Ṩ-`yH��Q�F�)P$�C�_���KX/�r��jHMQl�y��݂�u>A��(T�r=j�0�{�](�.�QV��DG����,�y'�����>�п��]��
Oy5h@����~x2��͝�'�JO��Ta~���c�l��ʼ~t�-��\G�C�vo�K�T7gZD�j����M�Ґ�2��7����4N	��aG��IʟmM/>�n�j��q ������wX� c��L�����J�=]���o��|����3'���d�z���QL�+,��M���t��U�j�Ic����B��H��2�f^� #�	I]�X~DzH�s.����<0�,��U�n��XG6]�\%�5�8�2'�֬�F �k>,ob�)"uT�����"��;R �S=e��kf~�5R����h��%�GɪfZ���� O�1�e)��S�����it��n����Hu�|v�k��l��Xӛ�_]�v05CS�vqtam���=�a9���v�%�y��z�qM1_��~��� ��;b&��}������dT��#���àoyB�=�7�=ᣀ��'� ��qr���)W|]z8F���e����j#��ް��Nn߂�Uj��#��p�;��ON��p=nܫ�&�w����W�.�W�}��E��&f�b]���_g�ԫ�@��=�o&|���'��B����"��e���6���cJnd�J���I�/��y��&�?j�����;��.)���AF�!�	S�
%_�������u��91�↶��Q�]*�� \ �*�@c���;�+m���gN�G������
\� a��~��P��%���.9�}��%E���W�b�|�,m?#�S �.\vma]$x΅d�'r(/�����[r؂,�w������}��H�:��3b�	AF���j+>��T�o�v�$�.�D�B�}rX�ĥ7�S�n����9�t:_
�D�ΠÂ1Tg�\��'3��!$O�|��	���f�����I��Iy����w� �h�������!�rM3����|�K���w��Õ���V|�	�2-��G�_�a^��������V��Pw�;\�l�g�ǷbyԜ�p�o��V�u��������y�!���� �R+��ೕK��˳�sf�ܿn�'�;=��+|0�vX��LtD����e_g�m�z�%-$�k:b�� ;hb%�K�偉�ۀ��Q�j����uj,&�����LA�J�'q;"����E�F�PKa.�-��֓��y�={4ۑ��t�F��W0�[�B�/|X-b�V��{F�Q��J���fn3����_�*>�+^��axC\���}����CRl��"��Fc��䄎��JȮ����b/~]8���eNo�n}����Б�́�Tst	��[�3����.��,ޒ�2����h���f�>���AV�6����`�Z�'-GSl�,+�Qw�҆ץ�����k�?�R��&���Z��8�g��h�8��5��,����r;��cg�M�4#-u;����o���G�� ���� �;RlB�}��v{,��@���8w��S�l�d�[���f��.���F|��VP�>�qy{��E��^�-����,�N��n��L�5p>aw�)��4���9��$���,^6��O�E�N�I���_cjJ�F��G��(��C�w�a;�[c`?�h����`S��3ǹJ�x�����THw��z˒�7{�=��%�.���Y�q�mz�3�B!��g��U廒�u��ϊ���}��en��[�U�����]�;D9�;Gb�n6w
	?�냟���sc�n̏�O�i�f�p��]��Z^f�Pp?W�ؾ�{7�y������rl�_���,�it^2�[�ޝ�4ߚ���k ���г �[�T?|����� L��7��_��i!'Cy��l������'ɱ�;��݌6�K���r�4NÕd�-�����@<�u��\��	��54H�p����G���#P�� D�-  ��	�H�]�����!��>��k�nd���htt��3�����:�,|�������q?�V;�Ϙ����~���ʩ!���E���������CdiǊ���;?�\{�\��i�o�"r��U������x�r�]n�Rx6P{����ZåI�{��[Qp���?���֯��N��V��h��L@Y$��B6����@�*õ�-�6]����XL����|�~�� ���3E�v�.�髭53ҋN/:��V��4-�ʏۉ������dsc7v�
��Nz�z�dr1]��N�+���^!���Z�cN^2h�f��m���?�@[�sl�c�%���(��[;�����R�x��~���E(�OGZ�(���P���]��|`�����FvP,��"����Fv��k�X�<���?a2��to���C�Wq��SǄ�H6(ֿ������3�~!���W���z�O5t�%����a���N��v;�1����k�����&;~���\�C�����#(Vٺ���
�TK�����R��̴�^ydm��P��=�ݨ��Ii��DV4l���C(�-�A
��A+?{��q�׽� �f��c�|��m�Y)ӗ�*%7N��^8�qI&x>q`K9��S��M%��M�Ό�j��V��(�0���ۆ�N�1�����(%3�8sR �D����/�"%~>a̱�֒s�k -sv�2G�V��c$�
1���+K=·�9T_��&�\�9����6T~@��ɡC(����ڳY��w�o�D��S��{4���������W�	b�Lm�v�u�ا�O�cW����wp�t?�.�mxn"Oa�U݋Xf��� �*����X���7�^��� k5�!����J��Wf�j�C����F�rhZ��T�:a�`<�L�I�պ���rf���
Sݫ�5hJ�BuЉ|!�_���dnF[[�\��f��rʂo�ώĈ�X��|²Ud��K� ������yծ������1�ة�W"�!��wG��N�;-8N|H�e�(� �L�#�$�+4F`�_���Sj�� �Wƭ�p6�����+e�����O�C�n+\�
��Y�&׽#C�]��%�fWh�%I�?���]�x&��H�p#u��3E<�Tn�+���[9_���V.�.<��#�������2+lp'/Yu�;w[E���cNZ�v��M���T�~
��
�v��	�gu�ƕB���q�#��|��TrS�H�������iΟ;+��7rh>����f�?�����we�<H��ܳ7L^�o�vA7g��v�
oz��~�ȵ˧�ށI��M�dS+��+Z�^O2�ʔ/t�p>!R`"%���/	���K<���Vy�o�<ɦ��䱐����]ï'��8����y[���j*�o,Ň�̩�<�J�����J�
n�ӷ��#�;���0�"�b�f����`��Є����V�#�P�N��[�	��G'�H���� 噜0���-$6�R��+d��%]w9vG(��J ���'�v���V����)W��qQ���9�)�3��5u*�L���hE<��w(
��7�2}2 �qŜw�����si����(�C��V"�ɗ�S��N��U��υ�Z�q���#���T/6\M?p8���fi�/�w�q���g�}D�T�����ؼ���rj[�W�ȗ(a��U@alypNm8���v{ �c��1����讖��U[I��iS��K�x�wަCN�79����[�m�ǔ�_����멺?�a�^�k���X��R;���_hM+߾U��FV}sP
;e{�-�y��V#
h*T@yH����TX��a�*�,��cC��F��_�AgG�Mm~?�X>��n�z3\ ����}ƾ�]�v��#��-�y��6���o{�~�>=J�a<Y9��,�[��y�E��h{߀<I�1p�� ���Bc޽?n��dӐHgO�HՒѬۈ_�8��~��)/"�S�r���Jܽ���y����i��u<�	�,���<"0qB����$*� �F�P�AXc��j, �v���C/ǠbR����Hw>��ݤ*@�1����ue�	����+?_��_�d'X-5�l�ͱ����#c��7j�`��.�W��g���A�x�M���T�Y���#|�M�ߔ�����g�bY�>�����QC���(���~Y��v���z�
��w��g�a��w����ʖa\�\�#�׌���a�i����i�!*'擣/�e�rN�<�l�0Ӓ���R����F�/�b�~����C�UZ�F�kn����*X�Լ�l�"_������w�����_�E
��YԢ���>K<�7_doˋ��]��NRk�O�*h�U Dݕ ����A=����|v�;�PWɠ��ޕюa%3g��.KJN7�3/l^���n�]��"����u_Ԓ�(�W�b������b�0����o�[�fifh7V-�,L{w,P�0J��h��H���H��(K.^���?f�p<��b	�5s/Dͦ�fb�����vO����(j�Fخf�Ӥ���p�$R4/�n��\@-���Q��;g&��7�<'�c���(�K+f��?����`�{�!qƟ���z?�������I) ����6l9�yQ}�|��kaU�����Q@p6�W}�Q��2��Fо�y�o���d�4��n<1����ĩq��w�1Y�g�j�#�ۊ7��!�.�'W�"�A�XL�:v"���������cv�"�
���68p,p �S�F��A�m�
����kC��:HL�𤷒������ �g#�r��2u�G@��᯼/:?.f6�fD|�}���C�M߾��:����n4�֥���n%"L���&�{��;b[�����qJx.�zNPK��X��k\Ö<��	��*�p�N�;z��]��$�{A?t���L(O���H媸=M�ơ X��%�L�\@�!��X�3 9��^;�T�N����[&��E�`=���G��WYq�	��CK{�]�D ,t�r~譳��� ����4b=��.OU�.`�5q�v�,�j1t8lH$�P���H�3]�_*���t����&�{'Ğl�^KK�̀3J��m/$�������ph&�<�G���\�#Ӈ�cd���>�K!AV����K�)�3�����X�]����!���\��#O�24�t�X7�%ɕ���� ��4��,~Z��g�>�3�k���l�#�
��p{����F{����T�]�K������8WA����I� rA�Z;�H��K5�,��i�}�L�4d�=-�:�{G�������@�}y�/�ݻ)����D��|mhq������~&���H��ÿb��l:W8W�[���Т ��]
㖫�8��U������[g��pu��.>u].`X�Ј +�r�F"������a.@;���H{-�@�g�\�φ'%E���m��5�69�<�����]��	�0�B吨D)I$�ާ����LQ�l����|�6k�Y~�DD��k�Y��3I�<�I⥶�A�|�{e3ŢZ�D��l��W-g��J.aFG�;��;ّ�M�L��m3��i*��,�3,���.��+����|E���o�oW�b��Z���+���Ly|��rD�ƚQy��o�cX�E����"3'_�cW��7�<���Ǿ�ӂ�%�:Ipr���X5a���X�{����,�HW�<��x� ��g�6M�r�g]�����?#/�4҃#Ǻa������2�W�)K�̻r��'8� R�Yp�a�\�4ˡ�$p�����2?ҙ�%���͋nR��jL*�BŒ���GY�d�$���T�;�w�# ���!@��Smh�/7)���BĖ���B#��0�ߤq����\�K�yu�՛�ȴ�(:,�Bv�hC���U>�V6I����YL�� �uYP�T��+s-�������)󶤠�~�q����dl��Ԓ,.������
8~��ƭ�P�>�g�@��R�* QcES���5v�!���`��C��4��>e���(�X"�*�h/�*8�}�:E��\�5cx+�H��)
 ��i@��UA� 2  ����A9 ��������֣�j�>��R����wh�i���`H��c:�Ej����*�����8D��[h�7Q�a�Z��(�9����,@����1 N�����6�%�����k�`�Ja4�Pď��� ��{��������d������yRwz�a߿��ӥ�t��X�sB�dB8
�%���;�)���S���!@�	z?�5;��|�(�U�J1�;Ii�	^��[y)loɵ���M^� -�����@v�-X�V
��L\n��p~{N�<�/���#�=v�y Ρؤ�K)����-���W2�\weP_Q�c�[�y���-j�y&0'��[���� �g��(�;$L(M�'v� Υ���!�G� �js�p&���!��
���t02��r ��4�i- g�L�֭�l�_h8�.ݷΒd�5�z���Q�5"U��J��RLm���G1(e�m%�(u�OG�d�[JU@���e�<m� �=� 'Zvt�gqsJ�>KHs�����Y�	�dC���z���'����3�O&��ί�e�~B�/�GFu[<צ��H�Q���kHB��%��U(��p��@l�Ȩ�%�&�ӛJ���)�� �OG��&�!��^u��:�*HD�z9nLf���3�>ƨl�Az� �覗�T�N�S�F��,�qQ��2�m�	w��t�lR�)���9"|4GI_;�%k����.'���+�.5x=��/Hm�[�pgU�F����EH=Ȟ�}ٛ��z7�M�|�� �Tc%8� �>;�Z�5))�pl��}td�r�TS�� �"9�@�ck)�Ώ���Q;�	"ݐ�p8�Ԙ���=?$vq?H=]\O͎�����hPf��jǷ�fd��<�.�J������D9�2�����y��A��r6%7Մ�f����zL"��#H�g%��Mx�%��(?�c���?T�v]�1�@N�,IVX�n��,���&p���?����r:�&t��Q�d�q�dh�Y\l�q����WӀz������o��������}�Q��1V�d2}o��!a2��'mxrGy���ߖʬMo�L̄��=�:K�4��(E�9��Ğ��N �S�CfrR@勪���)
9���,!��:~���`�@39Q:��}���n��6�˷.���D�<�D���=�%�U
�����PI: Q�ܢ�A�u�tj+v����`8օ��������:��-Pn�Mp0
s�G�܀j��d�,U0��l�)�0���c����Y��V�i�`�~�r!28��w�1SC�;h��6�)�y�;��\s��#;�m�g@���9���r�=�Yp:��N?���dT��b:}������h��pP�(H�iSF�2��(�_`\ģ�=�å[[�}��`��"� ��$���(藬�_=#�\�V)SX�R�	��B+lQd�G\���H��b.� �T�� �ޢ�
D�4�Ī?^wL��h��GF)�,�%�p������2� �:]_ �m�7�lfa�̡���_�k�S�R�H�`��L٥������_`�N|��L[�zVye�i�<�W��o5-=��b�tH����k�(Di��啼 ߃xx#���q����c4�x T��� k'Ie|O�^�UD�(��.�+ �����m̥��X�����xD�}"�_P��s�H��5PtEP_nX�k��W2 \����r�.lϛ\�e�Z
���]�5F��6���W*�����Z=�Bs�����6���0��tY!JȨ=��)�&��,�5��gܶ�:]d���X,��&B���{�K�绛���)�h����aNK�?z#���o�=��,���uj�����o�_X����5n�f�:xo���*�c��a뜤�XJ� d/���%�X�4��	�*��s5}��SA��L����5�pn5��/tDV57�sMԽ�ǥ�@.\���c�َ��J�� [iyXg·�gQ X���m�¾���N��� � �Bu���щW�z�w�.�~�)�M�nQG=b�!`Ҥ �^���Q���MڛQ]
@��K��E�"���Yb�;Ӟ=E��K]��zԁ�ƅ ��K��&62�1��rr�4 �ś�+J D%j��ϢD ��{�t,L���Y��7(����]�T�Fm��Ji (wV|��Y6�Wʦ��G����aϐ����|��Kvm4^���0@&*ǃ;B�p�ӄ*���X8��*9� ���
:O�e�d[�?ݵ��}��k�fY���!鵇�W�p;+n���!i����_{T.����SJQ=Q�Hd,!�%�t�M���n�K �ϟ����=|����@���Xm�z�c�wf2�Q����������~��qWB�	��������|x�h���a��J�� ��45U,�-�י:�^)�tG���R��|�z��{#2=��>28R�j��d���Z)u�� �+���ǰ,ͯ��� ��6�o�ȹf�O�i�����p#.~��Rh���w=���]�����p�}v�^���z�('C4�c)j�c�J
w��Sb��[g��D��-�}\�����gy��gQ{`�����;s���`�a�x��<���r��dE�:է��{�`	��(��M���e����@ܮV�^t������%�l�`�+��s�-b�������5�_�ꟑM�^����VC�P�ԋb��rFL�}[_�m��yQ����v���r�k0����3��#��A0X���6�D�4�k_G��˪cj��@,L
�E"Mc\�E���'v��(-E)�ӗ�Т���6V�����>X���7�!;�$g�ڴ�դ+��H���6V�؃)��<N�2 �V�vFI&'T�����{9M	lc0h�qաc�^4�����U��m 
��N��ώ�`I �Z��T_��)Yq����H�dLCh�
J\J�0�ź��0p���g �3V���� D��f%)(2���u|� �>u$�e$��U6���><��I	J���ڂ��?��>b�	�H����\�ne���(�4n�%ȸ�7�dWIqXc��>x�ق��	&���m�K3m��K��{��>R&@�mQ�f��_L�j8t�X u��o���2�M�bip��*g	�lJ��Sp�W֣AE�M�xBrG�qz���~a;��'��LEi�
�-D.����%���	�P/�p��SYfVVMօ�Фp�&�(X��Fb���{?��qA_���̄��ÜVM���뵉}{]<�sƓ�V&*�1�tӺ>�\����d��
��`���lN�5^b����;(� }�U�*ń��yFcR�!��:ʤ��4������u�9������/=H7�`�g:�l����o�w��7�!�C� �e�[w�Jͽ����g4A�0Z]ӧC�CDș�@韂s};�j晒��
��9�
�ڢpC�����t҂�侯0 TK�tg��RJRt�ؖ�K����"wpZ���)g��X��@��Ő!�0H�g�Q0
�r?m����ʸ��3�e�/��~�~0o ��3!H�@� �� N��Cl-V�j�h��`����2D�Ӻ�6��~b���DӞ��f=Q��>�ā��`"W�Q1��GP����Q^A0ژ2$֏d���G���N��Kr~.R�v�QuR 61y@��l?��V϶���?t�ћLc�k��J6�Rj&[0t]o����LgW� h�q�<����A���&�X"��zE��q�S�Q�޹FH��&��;��=�\��+����Rz��Ȱ@��
��[��)k��r�~�Dg7�x�9Vt�z����51�'9�꼐�Cu��7c�]_7�}�dN��W�]��?d��b=�ũQ�&l 6��";��}�����V4�sw�qָFױ]"�4|�*a��A�l�[pH�]�n��K0v�&j�ޟ�d^W{�<���FEm��ٮ�k���;��&��������	�}���HAc@4��W�`��led�PR�4�Or��b�%V,�	6���)T՗���*n�لߵ�ּ.nĭ��<7`��of�+gtK�œ_��坥�	N�Dq2j6�Z$�r��"d�[q�<ߣt�2� M�?Chd(X�D�;��"�?2�a|��W��$��SZ�orӠ��4��(�U6�(�n,�P5=�G� �d������t">Cd>����E�^䞨�}��*�o�@5����Lʥ̆�l��M%���ސ���*���OsJl�u���`pE�D��/��?�||z����+�f����PPYx��E6�'��wq)a�l�fy���W7�.�<����B	�)���x�lUѹ��ͽd��o�H���DW/��;t���(�k�J)��ؙ؛�GP�G�2��s�h�r<r�g�cm��������oGP&g�-�ٷ��S��|<ϗ>�͕J�A����it�G��2�Lۗ��F�a&x�wk}/��y�	��GQ��g�?x^a�x��F��C�l��-W���~"ڋ����6���k�����m�@e�B�����f;�O
�G�:Af3��t�,�?�[�Y�6]������b�����ֺc�<�7t��0>Q_�.�|�]ae�,q��������t�_��,_��PRla#q7N�a�ѫyk�[���@ɲr�����HEu�)&��pƋ��hn�ΊrC�uB�/��C�.���a��Ɯ
�cAxQ�"����8�y�-�*ʫ��r9
^d&�5%:q��k0x���^\kgu�[��d ^ԖH�nO�Z���F��7�>`�uJ4r�~[�:�fsՋ�$�{�oX�#@����;��e+�x)�����]se;[��E�+�5���Qz���H������;S��a�LvT��57��nOd<��ܼQ�b��%�� ��
"D�����k�R���Y�����F�� ]�'�YD�D��,�m6Ox����Hp?�Q����{k��֗"�t��G@s �B���I�	 ��5�#&������K����Yt��5u� V~A)���.gK�j�}S&s�׽l�eO4�mt�("	|v��^��^>F{M��� ��#|"즨Η{��#O<�����M��~���_TrB�$yʱ>��5��O��i�5������r�c��Z�<պ�[W�v?gVͅ��f�3^Hb�V�!u���I�
�T��L8�T��y���/r*(؊�6PU!�x����<��j0�|>�;,D;d�[l�������H���WK��\|�������@��ȍ��F�jn ?$z׏/%
����-7I�L��U+|�Q���o��rޜQ��O��8��.��S�P��B�/ҷr͐"�dN�8�N��|:�ȣ�zx��;g������8�#I_����\|��og�(8f�N���ˬ��o�0��D�k�O6&��쟛�tn���z���sH������ u��A�!vԀ��5�B��&�D��h���O�Md��,�=g��讅�65k̖>�C��蚹��,�T�:����-(/(���/�ƾ�E����#&��2�����s���4��'�\<��2b��<�S� �<V*��n�HOs��c������q�N�
1�B������dƕm.g�˱<T��Y���	�����O���ȉ�v��SaW�*.�ԗOי�xP�EcO�{�s����Ub�~�pG��p.����������.Ts�1�Lj��qyJ��.�<��杌�+R��]���q�J����l�쵧M�j&���������	c Ԟ4I�s�������
����+���q�j^.��K�����6|�(��4*�ƘQE}�e�|-��0�j��:۬�e����1]�ʻn���}I��s[��М�]d�k���!�x�ϑ눲�W�\X�[WT�N[b����>oct0�(�)%�m�.1j��'��P�Y�j�;_�A��u1�0�z(�.&N�>���`ޘ*��L=u���]m5��4^�r �xf�v7�}�XVY@0�3<%������t�٫�_��a��7V���":�_�r�azn�T���U[�yS�ǡ��C��_�Dr\~J�58M>~�����WI!&��/Ov�^���a��U��S�_H��!/���{�=�V�����	��0��<�����R;�\���O�|��-fLo�ܨ� �:�䫸��P)���|7��)ð������>8��b�v�~`��z`J���B&-U����t�`�����ˋ
���ƈ��ù{@5�m��Q�.�� B�H=�J���5��{	�tA�t��Q�^�K���sO������H���Z;�{�Y�9�\x��`)8QTɰo��ދ��*�_PY��&4!+�-���KNaSy �[0Q�`=�!9���D�TY�������سn/n@+���������
�b�w.��4p�j�W�]吅$� ����Y��܄��RZ<%P�H�7�
���
�"�GV;.��f��k�Q)�\������"���^�s&8�!�@�,���k@����w _�en���R���B��{�yj���2�n>�����<��]�zHٯ�c�Z� M9AHCX70=p�LBCK?ŝ�xV:���^�PC[5�,�k���P�y@?L*����,0!�m��rk�
�T��BGX�|<�	��O/�j�3�qQ@���ߐ�#�8�L���_�/~��{O���e>jA\5^?EBi������,�ׯ��Ñi��]&�5|ߑ�v��q"mBI0t�9@��(��n0�5��_b+��('��O��@�P4�5S\k��(%it����8���=�c�1��B�N_����d�u3dдWe�@8�oB��34�(4�ӿ1�bo=�����[1�EÒS��q{�5��Q��<�E�6��@������T|��d�M4!�#!�1j��m��m��H��#�n�2ms�P�u�D�ϋ*cRslL������[�8P:��K�~W����B]k��efʜn����_�&�Tw][y�.��>�پ]��m���>�_�2�����Zvb^�.f�U�hD�4^磚��r�>���M�H>�g�n���r�xOO��˭�-c��J.ZB����cS�I!]8H�{��M{�g��h�����06t��dvK��BJ��ػ6��r4�/�����};ǁ�u��'�-˒����e�|��Uu(A��Џ�g]��ag��؃���ٚ,�}�����¡��]�[�A-<�0J�����7�
6+p�&=?L��7�H�ӻ��Q�3�A�dx*��s�lD�z#�	9R>�I��]��\����>O��Jvu5�P`��x�k��UgERA&Г����8�V�"�C]>��(��{��tY0K�qx�9�Njs�ڤơk^��y(<�:�
�s�anK��ˎ�j+����M;U���f��y/o:]�xaq����pg�i�jU�l_Ќ3L��L8T���.���A�!�{����I����H1�;�25+o�*RC�K�Pτ�C* Q��T[.�n��?��^�"�'�e�������3�ķn��T[�D{�+Kcc·4,�L1�R
砪Z%«�Ó\�z�>z�{Y�Ԏp~w���o5}#G.��ii݉��"rQ�w0�j����8Xe�y��6�	DD ����7N��+�+O}��5w\@+�%?�2hx-�\�D�e��m��p�h�Z^.�i/E��
7*���^6�~ܚ�W��#"�.6/��_|��&r������#߷
�dlk��r6��rd�1M���J��úg�]�����faW��ձ_5�f��Wi)��y��A(�pY�}�!1Nlv�3��Oh�J�J��eMeM��]���7u�7ci?��Vf�[�"\l�ӑ,h$	��fu�v�(�P�F�-�ͧA�d(��X�2� �+�l�L(Wթ���N�U^��O�o�t*u��@�(Q�b��P�0mR�mHw쬬���*0,Wǆ�>U._�wsE�W>��G:�j�P6�C"�{2Usq[m$����^�ψ- �c���u`-���0"������D�ldO���r9E��l>ii��y��ZKه՚*S�B�~���B"d��O���t��{%igm�?zW�oF48Њ_s+<�?�t�9�V���*��+��b�8-k��r��  ��8��"/WI'����RN"9��]�5p�-&f��g�^�'�Z��_%M�AL!>����7n
0�)� F��R�@������:f�y�Ea��c6�Ĩ{�m�~��c�Gw���$Mc�� v�4�u�����zWA� �-�!�Eޗ��OY����e��{:�?��-�^Rԃ�K9�q��|Em%朄s
�oƋʜ�Lfج@4�ᅁڼ���.������y��k+�4��I�?�Q���k�*��*���6�����H��5��a��`2�����Q��T�-:�ֲ�Sang(9n����A����H�T���v���o�:�7�:&ݰ":�1�U����n���������BG��;�{ả,z��Q���Q��N��uM��ߨ�����!��I�����j���z�?��k.IC�1q=����$�pTV�W��t2@�J�]�_�i���:��ʅ��\�`����xB�])G�nM�g� �r|�{�<� 4�?E��S-�p� ������դtiM}[F����w,.��n.��{�;�ǚ��(��o���
�	�
PǺ3�_�X�'���ԀckL߾J��5����u��P��~�)[ܣ!�ÐI�%�"��!͂X|�P�5�-犵�#�R_dŘ�Ŗ)�;�t�-`���qv�I���@b��Y���A�c:�`P>�`$K�\�.B�U�R�Ȳ�����uw��ATI�Ps�7ߣtr���|D2�(Q�c��?J��{�yHH�<���Ho[9�*ٯ�.��S�Qai'���Խ��X�8Dc-˒�l��mzNd7c���ϧF�[�����H�=����g�R�3q����DZᝯ�U�E�l��}�;BI��w���/��{�c�����M!R�@腀��5���I�����Ы���Hމ�ˏ>9C��bZ�wty	��wФʾ��R�~�r�N���b�7�=����R�E�^����.�=h�����΃�������-����{~��s�Ζo�5�:�'�P��������t�=�f��ۥH	�[J��*��[fZ}�5sn�{Dk�,D�p�:�=�Be�H��f�����{��O���6�n��w0�ȭxyi��>Я>�}��')���F2�;��Qt��KQZv<�Չy�p��?�������}�1�GiT�:���,�WK�����M����l�ۊ�WV�g5i9�N5��h�3pX�-A��K�%�9�H��C�O`o��w��Z�½���0-� ��Y�99w-�^�޻f ��ip�q7��n�1���9H�<�dwQaG6tk�VyM�Ű��i��yqt�Q5i�?bp_O�����elʈ��K�m�\���s�R�|`w��|��gC���y���j���-G�s�'��m$�V�o�㍎;�\�Ճ��3�RJ�ؤ�,/�GU7:$^�������-c>I�h�6P�(i�˺��8��N0�>�B�۔�6�!�}f��R������LQ�[��� �uK1ih�[![�֦��Pl�/^^��]�}�(���8�$:XԾ?̮.�/H^Wu��?�lF���F��ch�gl���O����P��uLl�⹊E?e~e��#`�]����.�T-���g0a�~;�UJ)�Q�q�O������*S�ć� U��ONQx�R���C��7�KU/�zt�U:d�q���ons�N��$ą�=-��U82�s�!��HN^�-�|�#��/�yT��C���,H�����|���b8ڷ�WS�,��*I��el�M�?c�����՟����{��Htָ]s�0_�ۊc8���UV�������x,�ǟ1ɏ��6�e����p�f�8i%i���_V���� ���麺�����*�P���>�ۖ,����F�U|��nTT�ϻV��,�<t��)j�B��������.(4�aMaiQ��{��)�Rs/����e���l��c~�{Nt���8�G�l泜\�]��p�J�p"GN!�9���uH�x�M*�r,zx�A���%E��*J~+��Z⚂����nّ&�1$�#
�H��B�2�Қ�o+ҭco�S�	m�k��%RƔ0��9����/�:�f�-�O4_�0�6;ʟ�~�L�*R�HE�r���r6~=����X������
����b^)���{��:�2�`n�-��԰���C�ʑd�_�D�=�՟��G��ݔa���'p�5萠y�jA��iy��Ė�C��~�&�{n���}Z��b�������b>�}�<\��KٛkE���&����ͧf&�����N�Th�d|-P`��3$��yic���y-�R�I�o.c�?)��a\b��:�����c�/�����P�ڷ�f+��i�*Wn
N f�,y"�6H\�.d9���ǉI.�.d��>�i��I�>�LE]�3���P���>	�s�������w�#�wqM��Щi�~)�I�]��F���}(m��aܴ��y+�H0��Ǆ���o�ݮt2�]�>˭F��O_�?�a��J{TNrG{��Qy�׀x��=���*�Ec����Ql�����|�A��J����kPa�����������L�N��ʢ8����9�A;��7�L/��2�UG�(��'�lP��f��A��F�Sgo��]�7;kA�J��J��d(�Z��f)q.��flgG"���޾GS_�ō>ue%�<xp-J����z�#쳎�_�}6C��VT�x@��^� �l����>ӫ�/��Y/J�-�˒�or�§�*��-�d�|��������h�B�&j��
S�RTH�1#V���Պ"��nƏ�vΖR��D:�'^�K ����ڵ�d>�!'��
�Mc߅��2��ȇO���:˶j��f�5QV��.��5.�݉�^����Q"L�RQ�U�<���qin�j�݇bF	ĭ9K(u�R�Šx����u�N�5 �"7�T�d.��ͮk�l�D����Ȇ����Z�i�;M���;��\���2�x}������Gt��Weh-�]��J��g�k����}�"�:�����$�-��W5^�M?���,���~]x��7t��v� ��|"�E1_��R�����fB/u�RdQ4O�h���^w���w�
��"�O� |��I���h�qL ���'�.���bJ�	��)3���L}��32��TUf3}��9N�O,$�)���(��X�s�o������\��h{�@���1�x���{C�J)4�b7��<[�$d�����C�*��Ƙl�����BHnW���v��Q=t�&�c|�}M���R��Q٣Ob(n��Pq�Gq�.� �`�N"ӘƋo�"n��s֢_����b�dy��6y��ԤR-=G]��2Q��4)���B�r���V�EC33�ʙXg'���iP�yIMrޖ-^����8���7��Q�zm����2�M���G���[w�R���J/U�VV���
�e9�7���/6}�Բ��m�f���7�6�<��-�k�fAB��B��)**�f],F�D^:��2�	�õE,����%���ܿ�m��2���c�FtUfրw�c (�]Y����[3.�%���h�qG@�ɱU�ܦǟLP�ב��Z}��W��dݏQ�`Oh$��3_qjB|:�Tp�^I���F�N��+�f��XvP�읈ƈ	FG_"*{���0�><�L�-�� EF�Q�<12 ��q�?�2��"OW]A�S5�]��z����X�
tG"=g���޾S`_��9$��)��qҧ�F��Y>����u��S�Kۂ�PY�|:��5 K�ݚ�~�
+f`w�+ئź#�5|��>4:��<�՚���V|)�i�݀�1Jj>%ٜ;5E�5� �~.M�O>�����$�d�Dͪ���V��(M��콣�/�c�1v~wx�O���{ݠ'�fv��lQ��%%J�E��֍�A7W;�x%�33�%�@�k{�3�^�L�tp��fu�5'B^�ӨנmE�B�-)%�%����9���ϔ���1v�#��=�!�Z�G����淀�S���鵧�
 x�^�� ���h���#<UG*]�,�T�3cu�r��������~t��%M�xoU�8�M�����r�����������0�mD��������W2�Te;�~Ү�A�{lzW�����߳=��a�R)�q��;�5��(O$X�
6�Dl��P��dFd�o�PJ��X
��M͆-�<NH�5m#��S��B|�%�ܢ#��b��Ԍ��K�`�h�Vl'w-
���Cay.��|�B�L��9�Z�˅�v����w4L>͋���l�	ac��R�6�3�U�Hwq]D���0�6�"��0��9pw*}x��V'�8�_%<���Ż��t���W���3��q�]X-�t�#�.U�F;�ܺ��U5��������ٶ�����u����ܵ�I��|M���晸t���G�i�q$�MP|ϴ�MT�#�Y��}#��`��%�q��>�Z�w`��(*ʲI~�������ȼ�e��Z�-���a�|������Č�����d���Sa��\�7oʒٛ&"n��{;X�A�+ύ?�_Z�Z�8|;�/���\������UEǽP+k�W(�Ӊ��̓�m�6;B�ҦC�@�iw
��,S_��9"sa��Tn���~�p�O���S'���>�(_�/d$��ɣo�:xw똴�H��&��_�b.�����Ik[2�N?2�{~<���f���|��i`��+�	o��OK�6���ָq8�2V����V���#O�:��V�+�����r�;.pK��K,�*�c3D5[���2T3)��b���|��˞�B�?��X��?`�;u�]��'9�Y6Ř!4Z	��`�S��M�ψ��k��+����SwA��*��X���C��W+�����uT^6����ט�l^;s��H���̪�d(��Q-�|�G��b"J��Ec[[:J�b��ʉ��o?u�R�a�̱j����� ��|�����k��K����"�4�N�c���'Z�Q�K���͞ͅn&�� ]a�����7���N�MDŮ��_�9�9�Cl���Xi�	��7�61�h�z2�Q������tA9E�we�?t�`rm��y9��(���Y�H�h�O	��vu�.��;�%������f�Y`a�������?�'�M�HM�D�/���i6�T���#�J��7W<�M!�(�6�1�5�c��K|i������g��&�u?�gV�=��Y��Z!`2�O��V����M�e�c�#���>��>3�$��k���*�9<$�N�B4� �k��v`��5 ���yhm���pn��� '����}���D`&e�s������m�SgQP��"8gT���nL��uE�rbom��s��}�a?�pS���W?յ�;��^���	�"$�È�!���7ʕ�s�֏jG���CL�v���]�_~�"i���U����iM�,�mb�j��TE����m�U1����m[��'4�$�Q�c+�ۋ��t��鬜�[H�PſPK���%_K��+uĢ0X�����=1e��qX�ȖD`"�DI����59�t)_W��kV�h�8�}�c��~S�̈́��e�J��������櫩=9&�qh��T6ud�!/�����@��WX��;t1�(��ji����p�:�N&G���@�;6�S Je+���Y���o;�Ȃ
 �1�_�[������*@���b���ޙ_�i>�bC��_l�r�M%N����[���لi۪f������O�����������A`�ׇ���Q�V5\9��_�5��ǡ{W��e�I>ǇAy>����Sm�;�s١���J�b����X�;�����48y7��|�����<�!O��k W�GTFm��jy�}�B_�Y�.�3�#ٛ
~\�
Z'���;�+]6�+]�H���c�=��h��To��.B�"	���p����B���G��[�����j3�>��3��j��=~-F&���,H�P�~)�N�X�>1��"�������Э��C��v3stt�T���o�'��hӏ����9����� �Yd�J�P�c
j7D#�I�K�>��'ԱB��|��kx��ƕKnN�)Ԟ�>٠�\nR`��	X �l&�Wl��r�����E9\m�z$��H
�5���g�z'���( �����X#_Z���#����k�l��>J�1@�w��&$��O���D����5�R&�'�2O7Q�$dN�F	_	p#�֘.%�����h��,u3
CW�������h?��'W�i�u`
�4�VR�s������ !�����Z;Өemq�;��\������&ʜ�v�L�P����gX���<�r��E�`�n�^�E���y�0d)zTe��`�7�s�\�_��o���-7�km�J��@^0��wnE?t���[p�:Z���1�eq��J��^H�V5�x�*xV���sg���sd��5Wǅo9�,���uҧ��n~�Y�ơLj����(eo�f>�>�s����C��b�q��/rA��,����%�WAz}�����Z�ZI����m'��d JoH��,�9�r������Ir���H��J5ePEC�/O磻{�U�Fo��5����d��=����eދ"{n��0r��4s�]P7�r�N��|b��N��ж���ցj����_C=��ƃ*P=����{ma30�~�|�g�'�P���~K$����Ji���L׼A�Eu�S���7�O�ר3�vp���|Q��3t(�ji)DW��6K���&�n,Գ}�w�<S<ww����Y>��t�亙 ����(\�Q:#J���05��f��{>�'������&r��)>�&`Na�ﳼ jȣ�o�Æb'�?<L�7DM����X����|�ԓ��F�f,%����5�[V�����@��L�g^.���\��b��,&��ȓ�
���8U[����ޕUmp�`mW`dV�n���F��DZ����<M��r��_Љ�5|b�`����+�����_��m�ȧTV,v�bb����>9�>i� ��N�%�%�rTf��V�7K�7�C�<#�{"c�t,{�>h��T��t�����ȥ!�s��|�}�p�m��1\�c}?"��d��`��gB�釃Ǧ����FS����.���[�g=-S�EGQ.���WU�#��`>��%YM��%:(��N�5�H�H>`�]^��LMo��~�݇�nD���+e�o}�K*:�΄�n�N촏��#,�{"0�l��X���ٻ�z���R
��)��=�߼\ b&������$7C":��4�|R��A��J�b�ap�*׫Sp�IX*�5m9-�f[�dD+A>D����x�1�[�	]Z\@�[�X���	$�,e�,�©��G�JĀ�PY�!�wfZ�ڽ%Ozx
��"���B�{�B��<���p�V��~�t�Z�E�>�2��G���]a{I*M�W̊�j�:&{��TX�u�d�G�߸Ռ��YZ-�$�ꬍE�Ui�����i�i��iF���٩���jn�*=Q�*�k�����Ԛ��w�U3 	�Q��� �Q�)��!J�m��:`�'�7���괁���ږT�}ne�0��I`�������=�8��?����8�����av$;�.A&j��ٳ4x|�Үڐǟ��ո��p�l���Ğe���'ͼ��ռ��v�n_{�����-u�B���"I����Z��ȣ�{�+��+��ӑs�w#�;9�f&8Ր��c?�x���ܕe�n*���>���P ]��V\�s����#	]���-A�b��ق�Y���o���� ��A(~$�X�E>��"��V��Y�Ԃ��bo��x�6o�2���:Q�.��Y�Y1}���oI��Z��!p�)���g����R������w�v,�ͺ"F��AEb�K���@6^7�N�d���@��Ҝ{cQ=�'�i3�^�嚱t�K��������V��o�C2n�F���DX����Ej����N6
��~��l�����7�>^��WK[VW���k���x{��ت�G*�5`�6��l�{�C�����~�ި���I�V	����н%��k@R:�|C�7��BC��0�潩�t;�_s�+�ɞ��*���<�pmʷ�*�8�Y��|s���~�V�ɪ�{|H,��G0�T��,H�/ו�N�Ǟ�)U��!��*X�I��6u����{�/�sʛs_�H?�]��C"��g7�yҠ���	�v�����ɉ^gms��(�Y'[��`tK{�p��ǋ��������L@ �뎺���B󀟛�FD��>��\�+�3:��S�p�A����l�߂~���5��)���,�i&0����M��٫ު��[��,r�]���Ҕd�39����S6��_��M]tc$Kķm�V�f'���Oa�N��uZID��Ѕ$v�cR%�$S�dơ4;/S������{��M����|Sg��Z�Pc���yߴ̘q&N�%����7��#J�5`�����-!�)��+ݕlO>������vO�iJ &�m���x��Y�A][MGt��~�C9�f�'-��ӦJ�N̶��dJ�8�T�T��y-fIax` �1�����=���G���Z?�_�w�=�� ��y6`l�1v_ax�Hk����̘:�z��5$x��hUn�n�sv���Zam1<9����ˎ����{�]�����_�ƵO�x�%~U2,��à���ꠉZ�S�o�V[�����R��_�jAo��{�3!d�ZL�h�(C`%����ۙ=�� �f��C7HT6x��ֺ�XejTT�U�S��h��,���V�˴�M��DGǔ�����2�1�v��O�4>;��K�*�w'Һ�l4�;q�AE�Z"0�8h�j���: ��� �x�R%����&��S��5@�E#�*?�sJ�C[9�='�͇�~|����<�if�4ɩ�/��7�S��(���fS:U�s���
�Ӗ>ܝ�C���HS<�g�sDq�@G_�L�!㤆���m�~�=ԡ��	��̍r5~�V鈳��Q��G�l�V���g�Sj`�s]��-��`]�1�%�}�My�;��Z��g+�w����O���S3� ��G=&����|M|�����{)�g,�j���|+�)��0cf����%��	чaWYW�����,_��&E�W� �����$�]��HXSp6I�܌�t�,�Z^����17Q�d83R�d7���
���,�'�X�,�w�V&5$�L|6Ve�]v�$�
tW��� �ߒ:(���2S�D/�Y�.2��b�Uօ~"�5�s3�p'�l�M L�Z�pV����Էy�<��R1abG9�(��t>A��Ɠ&V�/%8�+������ĔѪ����4&�j�&

������mS;���͏��e�թ�����4"�ec�K"s�_�y����1R���jo�[��;� �s�w�k|׻<��E���U���J�� ��QQ=V̋2I*�^M3��M�+0<�a��#c�g椴ʺ�����DM���-Oxd��\�_O��s�k�tv���X�s5d@$ؿcuR@^D�V��?T�Ybs�L�;�'+�H����4���J�scQ�Y�16��n�i"�R��p����;c,k��{Е��v�]E9e�me^2�k���궇�ެܲ�˼��'ix{օ�X�����D� "��bV7��5�_�9[7��'O@!o��S�ɹ���!"ߧ�k>�D�,���Q�qJ>U�\yN���՟��|K��0����h�%��)� %�)�'�L�}>t��V��".\wa�3�ӳ[�Y�{�Ks�}�"�y�%ǥ�=ʐwȫBb�Χ���qo�U¥сUS�٘�v=��M�/eBߊ���D��Dit��*�1$�R8�@j���J!��cʒ���8�m[���r�|�w:Մ���d�Z?
��\��I��D��'�� KI���vO� �#�
����!d�,��o&:����&$ru��M�q�pOF�eF1������DW�.�_&�'x���?�v��0b}�����f���M)�7jSk�M5�V�z��@U��Q��k���G�e��5��
lA���+/�����.(C"�Gqz5�4��.Gl+����_��� 7�d��Ǧ3;��w~��W�n�9��K��{��˾�V�I��?\�`��t�cG1IT��io!��v:$z\���p��&x�[H�fd�э|?�q+g#h� �c;�)��|����o��fj_f���[�nQ������&>S�_/�۳ܻ"8g��b#7�}��W�`�I1�>(�Y��M)��x��)�rH����z��6�o;��r�����:��E����]N� w���qڌ�A��wwTt]�-���D$!5����y�<��$�ѪP�O�E��j�n�i]�cE,�0��Z�=�<���=)�,V���l�At�QR������͚�K{�݅���9�w,~g������{%*'aG�jt�q;��R�����lt�K�_�]5!�aŃ���Y^6�>H��ք��M��ǩ���6��0�^�h͔���'S�ށ����|��x-0�۠��v��ձ9�āX4f_������x�.:G���T�R;&�;b��Q�ko������=$�}�$��������nlX��^�� ��9�Ľ��<����P?�n�[t�i$�Qx��S"�"	_�|©�̗sZ�\��f�;���$�+�s_r�?����g��+�� � �(H:�)��6e�`^���"��]�<��'#q8�A�z0��7�PEp��~m��� v�e��FOy�0Z�?�-V����&�؂�\���
�A���_ ��"��?C���w��MfYk0.I�qH��\1/z�z=��-��[�9ܺq���n�,4���C'��p[�O�9��W���;x����qT�f���d������F��Zg���]��0��A@s�Za�߸P�.�-��[��9�9^]W��A�-�2�27�(�a�*��OKM��2��M�IA&�Ba��.�JJ @�h~7l�U<�:9.�DL@(�q��Z��,�ynL������� ;k�w�[LDkqWB��g�p:�=RZtT��	,%+V�l��r	�����s����S�l]����I*�d�?�q �$9�C
��>ܨ��ll1],bY+���Kl$��[Q�`�f���<-�#>ۘ���VN�<:Oz����:�q�G���p����oj_�����>:<��d6T�8�҅W�xa�69��@�o��)*�D�����vW�\I��
%�D��PWB8a��b���ƒ�~���]hX`�&�N�c�'c�!JR5K�� ���x$������\�i<�T�+@��OF�"�i�
P�9���%���T��l�-��3r����V覺0�X�@���'L;����%��ӕ $�H�.��y2����ǋ+�[I�kz�3ղ�a���O��Y)���Q
(�A��PcU,�g�o�;��}�;/����1hC������{�R��� ����Z{Na>�V�c��W�߈:�Mܪ˵���`&1}�u���m�x�`*U�
{�آ�B�,ٞ����9^��-�@j��^��-=�_l���M��RR�����5�n��l��j(�=#�"j������ߦL��5���(v�����5Go/2>����h�9�Ӷl�r<���b�#/?�ҁ���W裏z1�H��9�ٳ�W��N�F��܂�����#N��M�43����e| ��^�o����[�#:�6��OG������_���^*�*&@�c�cX��W��訳�ù�S����.03���Y�[YD�酊^1t�iȶ�b��g���y���3�˚o����֛V�e��Nj��tt�9F?Hx�������\�0��O�s..'ɋ���Y���.��?	�Kz�t�X������L}�M&�����\ML���2�5��3�k ��`�w��R�/&��i����v����w���b�V�E#{l��a ���t����ɥc�]K����p�5����ʈƽ!��h�W�W+�Gi̽�S��
>�Aq���l	93�׈�Xg�4�he�G�4_	�:3�v��+��8e-��}���"���R#��Ŏ�,����@2K0Y���v0��Y}m�<LNm��p��4��#F�URR�JYi�lp�o*��n�~'���W���2g%Ř[��h�|H���Qi���ʌ����#� �W�X�+����[w�źT.	��jAZ��	5fT�-v�Y�>�
�UӸ�]o�4e�˗;ˇ/������|l��^�',쌼rFj@Y�=BX�_t��83a)��������,�QÛ?�eY[lQ�3��_��?�O�c�i�����wzgcF�fp���l�N�3F
��9���&N
;0n�A�G�/m����k�� ��}���k�t���
�څ��T[Ⱦ�@H�k�Qj�4/9��T��\0m���
��6ǐg-a`�A�Ui���e��ֈk���oj[Ӎ�E��Ecj����w�g]�Q�� "�P�����Vv�=׻|���n��fXr���-d�
�M���fχ��^]N��|�$�� A��5Ĩ��R����_|KG:�<�(O׿�1��!������	;e�*j����S0#aE&|5�{Q�]�����&�̴%���ip��xU*)��9�V�-�+t����ov�R}��~������)8�В��ʱ� %'[Fj�oV�i�b�M ��PA	�5�m��
n�Ŕ���Oط���˸��hH�ldH�A}z�e�G�˔fG_§��D���O�9-�H��0�ؠD�Ḡ�f��](M(���s�[2I2�k�v��` ��ە���4�۟���#���i��ʳ��%����.Jw5I5�a��5��\s�gA�������,e�;m�+t���4eA�>뎏�_{�ᶂ��2}�����|��	s�hr{��V��ݗ@`|Zs"�Y�a�-�a�AEXf�`H������g��� =���Ȗ<��~n�3�wH���f(��i�ŲR�a��5��}`Fv�_m�� ��j��n������i�KN�����I�8�bQ��\�:�-b�+3J�uId5�+��{/����&[�`�52���BRW5\����.x�*$�7�����m�sq�8=׷�Ӄ<�aKy����(eb��Q����mK�|�(�.O��	+�^m&U �>�}���ѿk��ە��ɋsə%���}`=���� 	���3�~9�Qm]��nH�\)��J4����|�N�?ޤ�����xTy���w��5op�u� �]�"�a�S�9]!]���h������R���'����Jw�b��]V'�W3O�y=�ϑp��~���$23����
qP`�N�C���Ts�|�{a��a�ž�������	o���P�*�����1�-{���uY��9���������?&�{���*�C�|=ܓ��X�X��h�M�u��
=zw�^�&}���b������[�}�b+�v��crS�d|(Nf�.�b��2)�.�Zk����nd�I�o�}L౮|~|��xa�����>��'^a+�d���)���F��o�M�Gx�L���gA^�a�1��a]��W��'D�̜\��Udc�*��1ɛ�
Z{�V~U��d����|����Ͳ\��KTZ(fCt�z;H��x�_�i9�w�z;�}Hv���$�>�"x%� ����Ւ\���ʇ\s��Ec��ԛx:R	�F44W,�8�-�_=�)��T�M����)CHOU��}��.�,�0�;�T�s��(\�GcR��<�3x(f�-|�y17h�-�c�9���vJ�u#x#k��7I^�D;�^����������oap���(�9�(�m������qo��s�$-p������3�(k�bA�R�4��� ��5���߯f�����!�gL����A�ٸ�^ �n���͛��LS�1Wԓ��G�!�YU��_3��hho7���=�*�>\3I�(;
��|M�%iv�;��g�LVl�5`�g�`���K�j����W�O��2�Pni����Mƫ>�r� �#3o�櫜r'y���,��])�Ed����Y�ڥֹ:��h"}�"�U+Iq_��]����'?���+�0'!���~�nX��K1�_�Mz�f{�?vh����	�Y��;Tg�=��-ԛ~!�D�s�k�?��k���v��ݔ�_b�S�b����1�YCV~����fEg�߷�P�'ďA7}�އ��/����o����i�s��u��E"�H��ҭ���-tגX�\=��sk���('e:�D�n)�JYM��!(r��	|z�����;:����"��r�� �!f�H�9�Lv��
�HTP�j��IX�xĜ@^�b4�pÛ�b�|�sF�̬��;�ū�; ��{�b���_�u��Eݡy��28_z��T�*����i閔a�H O]��L��%�fұ�sZ���:�̋��Q*��+-�����0kw+:��A-�G��gr�:�ܺ�mV�Y*�F���{B۷�޳��&J��5K�̕E��˧)��.l�#/Fю��q�\^�K�;�������
����N�o��!����-�7��������g!��ҟ�h1��}v�b��b	>]ƿ�9x��:n764O��{"�������2,���{�(߯}t@�[�����i�N)�;����VT�;��nE�<�'�������9k���Z��<�}?̽�����|�Öo"�豂QW�p�����+��n��3F���JB�����4�s� #0����hf9;�טm�~\�u7yW��5i��%_��G�}quhUe����w�&�CŇ,�M��f'ī�"�*19��C1ã�t�ʔ�^��i�7a�V�1��w�U�C���)=����u��6���(Lj����h����)��U��EY1<����.%�(A܂(\1��걐ҳ��E�����\6��'f�Ӕ' ��A����^��(\��)<� �O*�N��tں:��{���{]��P���I�Q����sy��4�n�~AU����ra#���OU��e���J?���K{Ӫ��:	v(XZ�(b1��p��K`9�d�N{����S�ҩ�E����mB0�Z7hgۈ3��݌1��S�dVzp�X�n5���8������N�2V`m%!y��c$�hM�p��X3�D�]���8kϽ]g��A%��'ٯ�.07�5�v����N��]���H��G���P]^#��0�q���U9��Yg,��y����)%�߸�=eI�+���2T��K�9��g�@��[�I�L�@�Ss�.n�L
���_�����]Q��H����O�2u�oN%j���K�
�TU�Y���vc�?:n2��~���	�8e[,��j�;�c��xy�F	�ó���[ ��?lv�z��: ]bG�C���ؑu� D��@���m%f��	�����v��bN�`lCA�fV�k���GJ��L:/�P~9Kh/\%��h���GJ:I.�S�)S�` ��n\�A�;h��0ϫ�cݰ���rܻ��Y��i�_p�	$q�޿�;�(Y�N���B�����8���B���dͬ�[@�鳈"�wn���qE�'s��qn1ŧ*���CU����C��I�\�0b��fbj7U�:x8C�������X�`NB�x���G֗l�Ͳ�dȧ��x�p��2{�)�"<��ь�(�)������5�嵢N*���N\�G��хܫ�Jo�tD
����߬��9�3�׾/H9P����q����D�[�-`eI�����K��%øc�I�m���]u��G6�=J}x������${��.Y�l�|���km�/� ��)�-�_��������0�|�Tx���5VV3�5zI���"����H�i.{�5�=�3dEokb�I�&��c��XTV:y��y}bI�29Q�n��*��C�(�V��υC��UϒlXHѣ��ȧ=�����j]�C4��S�'sDy���B����W��|.#f��(������p�_��cۖ�]A�(Y(���l�}rb�uxXۦ��2rV�;t�_^�����_r�W�L���9�Ϧy�X����y����HA-Wܷ�/�hZ���۾���3���0>�ؔY�kበW��s�d㯬�����Tvdf���^��)�\��~�%;��G0�=qg(����*�l�s�T|pc)}&R�	JC'�����?g�n�	��Ƥ���_�|{oh����S�j���f���Y�e�w�=��wZ���-Y����|���:��������oT�~��=�������[�X�<�L�	�9r�_R=��)�6�Ѷ���B�|Gə{��*n"y�!�^J�IYb�|���Xf?T�К�/~��W�L���J��#|��9ନ�dE$nFDnh4�i�v��1�V^OP[���7Ά��z��*ks�gX���=�h5�P��Fݛ(��f��J:���s�"��t#49yI���c{H��I�q����+DybEwX4��ڳ'�[TI):��dV�e�[0{tm�j*��b�d�or���L�8ś)��w�L�v��T�1�Q4'P"��u?�Vp�k
���0�gg{4�w,<|��U�O� 	�T��~F QM��u�k��|�E�)��8̛h���(.�4��֘���&��]M��␃��X��8���dX zz	%�]�4OU�ʪ$[z0�A�P�:�{am�3�����"2���XS]s�1�sk���d{#-'��pc	����ð\v�����Dm^�˺V���v�g�<=Ib��	dE��ת�4�DE�������� AbA���� iST�ڱ�}/����J4�k�Dji�UTLU����d�*lFESOY��p�Mp8奠h?����z}�iC&�%"V*��J��L@�dE�V�i�R�tG7o�kBuv������e1��Vp���;
1�`&��m�2~�XeO<ǒ�f�Nߘ�R��O��;���ءf� �!Ef���,��T��w�F���W�fwC�4�X�&�؅R5Ľg5�Gs��N��s; ������3Q��\=�"z��cώʅ�ٸ�.�c\ ���HH���  8 �\>W<|j^m��RZn	��:fH��k	��5�u͉���-����?a��VO߱�=�;L��5�T����=vHr�"7E�,߄��:����#����"�{�h�<��=���
��U=� ���͌���\"|X�̫s�7d
mi�U��y/���*/�?�N�w�sy�3,2��/6�f�4������Z���j�S��� "c�����p�S�f���!�m�t�U�;���jf������-��;hC�\ѐb�I�aQ����q|E&3y"�Q�D
N�D��\^�T���Mf���<T�|���K8C"%�v�K.�)J��6~�+�7*6��̌��>\�
g0�	�b�7�d?���@�%)�{�C�?,�F�إ��\�+x���hi[(JF���0-$�������=�/u�n�&�/��6�3ا3[�}��� j��V���n���b�1���M�@��"�-9<h>g4�gf'���G#�Ⱥ�Γ���X�M1A���*~<<q]Ƅ�-� �*��eK�t��&d��A �+��6�Z$��[:ݏ�K�o<�G��P�Y��=�b��<Ud����/\��]���<�Ab	���[�T}i�$m�E�w5/��ƿ^�ˇ&%�՟b',�Vq�h_A�m�����S��C8�lo��)(�?� C�v�$��~'��Ů���ėr�8��}�Aiѧ�ćh�:�C�1&��Q�~����Zٷ�Vl�D�Q�H5�(��"p��ܜ���c�K��-*]�T�٥_ankB|d���Z�{T����*��{LR�����|��e0F��j�[&:9��s��󖢷 ��O[L�15�d����m�v��Ã�B��玪|o�`� �eYP:�'��&��T��$���6RQ c��}2���Jd#ϣ�I���(�kY��:�B�r���D����(���rY9�<TS�b��	��@�N�$��2W�_�jUS�Z����a�+�*kL�j<�H�y���,�H��?K7u���!��x}�g����5�>�SH��l7J�i��؅%i��`�rc���&����ȱtgfW�Ɖ�Q�y`}(ʰ�Pf��Q���
o��g/)KRŏV��GO���S��BlcW����3eה�F�U������R��#��ym�'(@3tY¹{�>�tW#x�)!	��8|��N�����@�NN
��q��I$��V���=�'zzznzO؟{�PR�V��>b�R.hW^^р��%�Ǔ7ŏ�հ$��|ê�.PG �3&��?�.�0�͆�G�+L9|��}�_�uB����)d���h�dENY��J m�PR����$��e.}����)=F��։<�ű:�HQY�߶]&@A�/S����u��Qu�VW]�\���� "�U���ô��`����%�����.�i�O���Y���	����J޾�JƜ��ѷ��^����"r����q�a�.��%V�!��S�˱SW���1�q=fٗ�X1�"[�ҹ��'a6c3k�/�rش�\�n�&�Y�$��2l�$e�_�� ��ߤ~}pz��.�L�y{d���M�u��\ щ!�׋��{{�p˷���^��l�GSFP��=;F��Vs���ˍEr��jy D�q���Z젍�����=wX>{d/��1������`��.2�+�m7���]{�ɯW���Bᦊ��fj&��Z�*���M�_l�)�'D�C{]��ίn���T�6���8��6$X��/�a�i-�|P���ݫ_�(��Q����h�1���/��W�xZ���wd��jL5���&�c��b[Ӏ건��12�ͻ �<*������)�[��M�6�+4�2�^\�t��M]yQV�*s���[u�#���u8�ʆ�d?O4H�Q�觿�������K�9 ��C!8|E�oZ��ބ�i:u>�Kg�B����-�)Q^ؐ���0DMI[*P�
Y��U<��E$C��e>��E�V�\+�ʷ�I�W3�.�M#�lr�
�;�j�D͢�͢:�R#��k~6�A����'`�8UQ�$��!{����:x.�UdA��P\���+N��'�d.
��&lu�)�Ş&�Iߺ��mdү������q�*�|p��b^w�`Y�E�D�p�i3���	Y�5�ʶor���,�+��k;�=6-���jd�#���*����o���e��e�� {�ڿ �
��ﱫd���i���+�gV�s'O�]���jg��z���^�-��9����4U��
�<RCTj9�޾{�$��5�㷇?��<���������ogT)�:�A^�t���p���6�d<���*�V���ml'W͵W�7Y_T�2��;�O��ţ�@y�QqNCgGeE��3D)��'La�=�Q�98�ԇM@kOC@�ƫRUH���*9]�)w�kmٞ��H�;Շ�V�� �E�%������Dv����>�� �o2_��J�X��6�ٮ_8��t��-�V=�\
"������P�(���Px��d�Է.��
��P�6�K����/��a������`8�u�r '�.��Z�#�e ^}�Q���d���ši��IԱ\I���[���%��%�P�y��K�ܭn�/m��C��ҷ�k��{�Y*s������D��,���E	���wBv=�H�A��݋>�(�/���*Lbo�Rڟ�J��|mQ�O����,��P����H@�y�h�5Y/1SY�8C��h�6�L2yZ�"�uȁ���H����/��X�rf:��@DW���QW�J�>�'��k����PE�Nİ��B�ee�}6�O��*|T�P��r��c�x<�q��>�
���_vW✜���Z����,9?��_���=k�� �ѽ.wL���r/OQqD��%��s�e�<U�c+4�6���c��������t�4�u�x�s]o����+R��>�c�`3�;�4GO1k�89><8v�.����ܘ��G�l�Q�>�n'f��q-�N��%�<�iN�+ܼNt�C�(MN�lp3�����#%�<�]���#bE���R��[���g�j��%�AAu[�Sr�/�5������C� w��1ۣ����g+%T������3/�v{��<��=\_g��݁:X;��ڛ�u��>v5�D䐤��0���X�vQ��(���#��X���wJ�s"_EAv]�o�w���oE���/��̽�d��e*�d+����y15��8��Z��/��
AX+�g=�$�_�������3�^��|
�Ls�xq��ҏ�L-tТ���:��GN��`G���7��Y���s�k��ϐ}(q|�e�đs���ʚ^(��4�	�n���)w�ҋ�i�ߧ�Y|J$��"|V~�a�����R�H�jP�+ p�(�):A�ֲ�y�y��ʕWv$�l��v䅈�b�ɲ�k=tV{���0�̞��F\�����:��{�!�59��/�B�����M}K8g�m'�vhۋ�h�7������A�&?�����
9��c�{���uB�K~�9�,܃M�]�r�M�`�އ�X4d�/���V���������(�z"(�=�1坝�΋o��!F��I���z�Q��e�2�4 $�L�$��[����F�P͐�d�ݲ�Z���� �6��@P���i�TnR�sD��uhtV0�)ǾoL��E���,s��`�/$XV���e-v81�+�t��G�rB�m'2LOr4��t�WU����X>���7TZ�u�Y+ܡW)��E�F��I0�%�˃���D�	��[@���~߁R=�|]�jX|�/��{J�{$��9ev�{.�I�N/�S8uw�5�b(?��c?��/�����2ٝ�"�'|O��!��1����'O��7�x_�eŻ<��|�Q�%���YUVe���w��ʳ-��>��hJ�s6���M;n��*el&�d�X�n�i�G@N���O�-�肦L�s/�
�'x�� /ٺ�763�F��[��r�	��c�#mG\lה�����I1�c�{���nRʜ�bu�XX}h�}����=�#.}���?u��a�֬0�VJ��+a�:��ړ6(Y����MX��:X�#ļzZs�i�η��)�恒pH��Tt��zY`�hU^m�[uG���c}�x�Jux�0R�oQsS'���bn�>���_?��⇦O��{�0��k��T ���'t`(r���a��!,j*��}��ۿ�3F�#���4<8!a��P)�w��8�L�C����2���>D!\͊ޛjq|I��&ʫ���5g�v�ȁ'*�@]�AF�s�f�z���?�DASv4����raP��,<�Edմ�p }>Z:jU�x-��AQ��7gm��b�W��A؊E���:e
��͌)�Ǥ��睈�g떽6��=dp�9��}����[��?����l����1����%U֗7�k�-��d	i���Ka+J��e�,�\*`���4@�a�Hx��?��X�o_�}������µ���c���c���J�)���۸���4/j�Ҳ���0,<*����j�gz�c~V�r�ņ����F�B��"�D����F�ҦVU��\u3�c�s*v��R��z%���*Y�8sC��ș�o,��-��U�Y��M��O�4�,]�Z��#�n����Y%�Y��}�,l>�{ɦ+��@X�YY�^B�F�n��Z���*�C����V���~g��2�o�C� ������`�x��N�l�[q��,b;\��G������N��.�K􌾐�[�(�6�}�����?H�aI�������և�!���(H3ӛ��(���b�_l�~����#8T:�ם�wQ�/�Kp�(�>t5��o�^3�Au!d�pQ7����>~�߽�62s9�x%G��6`�s�|�������*"�˓V��*C��� �N����w�$��ZJA�5SN��(�۫r�^f5!L���x$8���)FP�ҏ�h�Dɚ���f���u`h�`ɔ!g$�~n��]}/�SK���}��M�>����;�ck�92+��˱[Ox;�-/c��&|3��m�r&��tų(lOh	dvs4h]8*���Z$�m4FK;��H�_$�b��Jq� M	��F�Z�P��ITz����@�"r�{o�\��62����%���NE߹�$��¹y�v6���rG�hhQ'��ֿJ�+LE>��j}ɏ�P�4��䉼<S,#���?*97QA�/(2�ԯ��mܶR膙e�|��NE��S�)�B�3�{�.U�?��s�a27D���
i����2���Nf��]K�`%�{#������_�֟j��8Ĕ�7��˫���g܅aE���p��Y�?Qww#��V��m��x�b��-�e����-`����-�[�Q��U�";_8����:{
m���n��#NB�ڠ��!0�w`jaF�x��A�4����J흕��>�����a��ֱB�3��Ί$E��ci���`���a��/'w�.�Ϥƻ��瓙->�;"���/�b3d��<rR�И=������$q��/t�@�婇p��J��C�T�i���&z�ʁh0W�Ɗ�ᮥc���Kl��E�	q�ml2�?v�#��va����>�7��o����6��5Ӂ�7�`� 9�5%�!�����:��Eio���/�?,-0�7�s��Pd�U��m��lF��t{|�w����A�Y���<!�� ��"��m��^�Kcp+��*���W��}JY�e�G�B��~w2(��#+Ǆ�XSbz�$��DFX)����A(�,�����n8Ɛ�e~m1A��N�.q��*F���e�����=�X#��6�΀���6�fr� �Z�~�C/� �7GԕW%N�+	���\ؐ~�使sAcK����2l�Ǽ���u���tNA,M|*Q�J�opX����[��`�O�5%��Z��S�Fj��^��ݢ�(��)���Y�2�l���u³^V WO��
.C��H6�M��5ɚ���s���`s�ȼҜ�Ws�R��iX���4�O(j�Jb��7j� vS����\/9��N\��Wz�YQ*υ"nQz�F�0f��	tU�� %(�|��y ]�*�����o�|�G����#=�>0˾���6|*��Aƴ�/3=�B����B�T�M���IWh����_�|��|L{0 g�r�@|�Vq�w�<3���*v��kyyEʟ���M����lڦO�Xب�L���82z4ͩ��X��sF��~���U���ـ��{�b�1bh��)F(�YpZ�v�����-�X�U�[�!���L�R�!{��QD�������y-��"ؐI����P#s/[�y���{�==n��_�q	k��:��|Xre�PG�O�[BW��P�r�N�0Z�һ��[��^m�L
O��}�^�3E_2�H\�a�v���(x��!�dE���*w�S6ݸ�*mI���	�g�܊��
[�eT��� �s�ӻ�+<�H�����$���QPX�{8%�)^��$N�.��%�p=�Z�i᥉�3�M�]B�,|��ݗ6���)W�U4�eƖ��~E�9:�xo�d�'ʻ-����Ւ�A���z����3��-\�n:�_4<'�9�F�nI��7��Z��}�`��C����4���`�8~���#&����Ԏir�/�g���UO�����+-P��ށ���ޭ�ä{g޶e�޾)9����_����q?=��n҂0���u�Z,HC��R���y����x�iXK��zb}��j�qr������cn0��K=�9~��f%�>�!>S�5gWw�P�'�6���e����R�a�%��T��#�g~��"T��i��Y}Z��$j]8 7Kvk�Sr��.����I�Q���.�(��N����1$:XkH�M��֞1��O	ð�֚e+f<~��Q7b�,�[P��X͕��5�-�j%��!b�����9�gAI&����鎊�$'���Y�C�Vű��?Hκ)�_�ҋo����R�r=6�c�1�����ߟPv���\�[hb�����68]p���M���n�\����� j��o��R-	�p����۽[�R��>����$z�Ύ���Vha|P��7��Qr��dB߾Uy�Kɰz�M`���R9둜q�7��Bp���e�8�+������M}�qkA-�PS��H�M��\O�֒���s�ˍF���_T��|C��R���цi�'��; ����B���e��k;"�ģt!�s`H&䲌]��W>�˃�)�%���W�3�y�rƤ�(Ya$�g��D�1 W Z� "�N^LG:T{nЫ���/�s�[q|��r :=�z8aq�u���oN�qX+�/y�b�x�r*t~�y�'�O�7�eC~j(��?B�Ȑ���soc!��hE�('a���,+���n3�������TǄ*�%�k����Y�؈m�]�ScNu�'��_1��idNp�#Z�o�d8�6G�޷��{��;�kM*D�� ���?wɳӿa7^��g�Pm��I�m�t��U��1�1���c_"��9��jG�=�z��R�z���������7���_�I]X�|϶���V���AFo[��Em\iL?R=0�������"[����4l��x�:�����dX-�̪�V��,�l)�����:t\>ߐ}�O���L%2u�)@~����ʑ��h������ nC�0e��0�:M!�_w�uQ��9�C��1���������>�m�%Z!t�9�$ә�2��7���zw�D������7�7�ȼ���e�-ZE��c���W����v�)H�Zk�6�R��`9�Li�i�&�n�ظD�$$�9�q/؈�Q���_����ʣ�i��;M�HH$��z��J��=��t,0=4<w���:���}y���6׷�=��>�AB��y���l03'K1�mr�R=�����ѽ	'�g��d��ޗ���J�®_#:l9��5�J7.R�x:l���R�Q��)9�	�vZm�<��x�f2� [+l�7���G�8
q~�le�usV[�Z��s�kR?��mM��C#�����'��%Uf0��m���u��9B�ơC��aM��x��?�E�߰FD �ZE�ڧvNEUjS��ɇ�b�Ё1 �]��Ic�Y�����s��q� �E"w��gM��=�O�ۍa�`�vEٞ��(�ڛ�P��*8���gL	�� ��ɩ�k����iK��A:4�PG��Zߦ`�W�:��p�5���]��ӥ�J[�gv�d�D6�����Kndخ������o�-H�q��mh|�v?1.LR�x����ǧ��=|kn,��Q���-q˺������������˩���f�s�eI�9��iԔƌm4��� �r��u0�A�Qʀ*�_���WƔV�'9�Z��(0}64���f��D�u$���(f��h��m@ @�CFC@Dx ��� ��O��8��<|�x�4ܼ�Z�n���h4uܥ�����1G����̯�x�Wp 8IxD3�M�A�|%�]�|��§2��GPt+�	_x=��<0�kY]m<�<ߐ��;������H-�Z_7��jwH�g;n"\��㚖X�ٰ��ڢ�zh�,!��:���!V��]��ZG������)�L�4�s���
| 6�A�)*D�Yr�x�f۝�{�y;��ݱ�du�aV%˔�n�N�cQ_W�\���PU2_*��r�H��Ț7`횰f(6m�#ʗ�SGh%�a*1@�	կ\p�L�wE\V�gM�a��o'�u\צI_���Q}���v�x�4a��?}�n��b�Ȁʚ(�T^�J�	���wȥ���Z�t�	?�ˍ���I�C���e�EA��>b�ƻ���"��O�����ɒ�,8�}����xx!�[��� s�q�!c��%؟=~�uQ{l�o���ه��Ӕ$�g�El�Z��iU�_IK�����\���:+�1"��<=D��$�+��������暄��"d��� A~K�xӛg��E}Z��,Y)]M�*�f�7�E�[4^٘I}r�y"�8���3w%ڨ���J�q*��˳KY:�qn�!Q��A,�L�$]m*+.(���P�8��[~��gX����xL#�8	7e���g�L3Eco�h_��0��3[�u*މl����8�Q9Z��|Xe W��rڙ�F�����K8�`���z/�R�^3���(3�G0�|���Py��z���v��.�-��ɸ(������Nq�Zx���9�xw�S?�����*����l����;o�x�����	��i����^��s���������h�+�}���&`�W�hs,h�cQ�|:�k�_�B2���� o�A��""ǋ&Z~R*��Q�5O&�yM�P���|D�h_�ʍ��"�'����/U�������p\:���#����i�$�e����I�̪vyPЪF�X-Ӱ�I)���2\������\+p�%�YJ|A;��M �)e	��1>��v�w��l�3z�����[�Ŏ7�,�L�Dކ!#G
�u����]H�H-ג@l���+^f��R�ĴxYy�«T5T��~cRRs=��3'�\|�n;[�}�J�i�	!�p�����*H�<��ls�w%�I������R5��M��{y6h$�.�Y�6l$=.y�=U|�s��yw4���@k0�g�v̚@�yF��2�Y�+��p��	\���].9���Y��y�_�/�#�{��{*P��x����Qrh�w78^�����y�q��$isMP�\�0���Y�5�ǭ�	��ى2�S�U,��S���ɠ�;�X4�]*���-� +��tx�ꫫ�2@��K,�JൢJM���Yv�|?t�f(񽒇�M{��7�x=L�"�c 6��k����w��Ѫ?���X|�
ڑ��������5�GY�3��i��0\G��.�-�٘�����u%����
��*�;���Ǘ���k�B�2��q�t�(��f�6���KI&<�d����f��#e��ڿ%З�h�%��B�h���n0�8EQ˽I+u����f��O��g��,��O��6��{X:�'4Ff�������7�������0QЕ&z�t�	�}D����*�	���λ�Pr�4����@L4^��#�T�3I�w$�������9a]�m�l\/���H��Jj�6Ny����7�����R���w�}�U�z��\c|$A��f(5V4f!z�%HՁ;��O� ��l�i^ɆPF�Z���Ր�mm��*뉩��5��F�T��s-
-�ș�AY����'��r�� Q^ą��Xwy�g���8������_�q�0��zM<,+=�4P~5
7Kg�C>B�i�w� 7i�=���8�Z�j��X*���$��� �������/��]���֖��d�(琖Z{8��{Qٔ�YyS̓�z��-�_DMN)�#bYB�~G �R��s��"�O��P%�yi4���,3����d�.m���&����w=i�ӧ�W�p
��2N���⩵~Th�C�Z'�"G@�bt�����^:�һ�I�Z$,4��<%���@�NW\�n�E�e�"�:ւ<�e0��_r��ۚ��l��y�f]8�p�d��g"E(�-�{r��mꗅC<�]�r���}�J�"�o䢓I���M<�"�DK�~\ǡ�����O��򙻷���ų��h1&+�;Y)֕�i��t�.���=��J��S�i�s+��"�­OyL�mP�V���Ng{2)�T=:똏 9-&�9���PP�\Ȅ,�,��.�d���ev1}�Z��g���Nr�;�DJFsp�G��Z�?n�T<<�ycI���l<]�ll��fP�9*��e��e�}�p̀R�b��@��B{6N�8�J�<eY��O�E�����jA�^1͆9h�t$����@�e ͺ�4{�k��u��`VL����pY���~J��>ZG*��ƛ̬�����T�%V�J�K@Ų�D�מ�����}X������[Qdߤ�i������7p㔳��o�Q����"RZ!��K�*1-��1J���ʨg��㕦���GH� ����Z�I��S�0��Ae�?O���M��<��A�U�Pzc�$T�@ŕ��HYB�j�/�����u�%2~d�>֤�Z��R�)��}���v�F�V�S�t�7�O��M���V��N��9�����XMq�b�&���2��T���p>S�܎�蛇G7+U4�c6(D���&}QD��H��5ʹ���jI(7����i�+�T����fy(�_%��/��~�_Mbଅ�L��֭�>��u�)�ԥ����.�"��a���>�Ġ��$}�A]�I��a?O��A�cB�)q�+�$g�����о�z�(O9+1K�5����v��}�i�������'��;�y�⭒��I�0�--�y������Y�I�Jf��`T3��`��!aʒ�P]��Y��>R�K��X|������!����Bj�Gx?ʰ늍�sg��2���Zg>�z@��5�Fכ<&�c����(��TbA���	$~�>�C7dP�hj���?��a�������=i@���^U�>��Q��E��₈����i-M�P6}<���P�4Qj�~ATSQ>��p'D��J�u��U���>	P$�U]ۇjzک[p�9�$J �n��N�D��2��,#��tzƈ ���ӖW��ET$����%��	�5t�JQ��>���u����r����.&��J�v��l��F%<�*��.���<Ra��&8e��؏Q;�H�2v�S��|Vs�����O���޻{��6}M����υ��"��_�A�&�2���O�ݡ��Q�,~˘mD�!m��P=��,��`=��7�ɴC�aۏ��I�,�=�-�E�hZ9�5*�Իν��p?4��|\���?vxv�٤����H�ʉ�2�	�Y�ma��5 Y�$�~��ݩx�j_���{M��m+<n��l�B!Ө��J I�Qb��y�3Ѭ�e����xP6�ꄽ��
R�$ּCVi�<)�=����)�G�<�E$�^y����]L��bz0$u��D���%�r,��i{Qwpb[�x��w�B�%T�puR��rF%�!0�J�u���R@�覱v����M����^�D�?9�2p����2���W=�i5�5n}/�<~m�`)���%��̀�e�~Z��p˒��o4�Y^���_K���v[��.+ T����6�y�E������'�ޡr��T���2�����J���W7�w�b��4����!�cԆ�%�/�R�^b$�LM_�u�7�B�P�ѻr:�`mTl�-�xn���]46\�@B�q��X���f%M����q�cs�Vgh�
��qΈ�gr�s̳��/��pΙ;Յ�M��pKp��
��p>��̏����.	���C��Wb����3=�B��0 �;�F	̓�㽁|V�ϻ��&>V�d���a`�.����s�JȐ}YOQX�v���SvPn�z��O�����8��v�F�t(��}�kun�A��Z�� �_X��R4f�(�M&�y��V�ߘ^b��L��̢м4p-?����Ly�iϚ�,�b]�$�c&p��i�����W ���&�/�|D�rT�T9h��Ϳ��3�����![��z7�h#&Y���B��0;�L0��c��q�SZ(Y��(�e�'Kd�˝�ȝ�b���[C�Q�_�6��Nm�銯��+���z��Et�����B��ltD�P�-r!FSԖ�O�Аuq}tE�?V�����v���a6Z��B�%�%�ŗ���f4wk�C-�'����:�G�PA8���k��(J�_`9$n0���׺�8u�u�l���)?�O��b0,���}Kx3{s�ᘺ�"�X��b�����"����Ym��o�h�}�t�H>p[�ʽ�e�y��F�'��h���׼~���a�'Zwn��g)���p��������7n{
8�,)+�"NM�~��Y�O>�HIe`��|�LCf��dk|�6�D���Vd�p�2TQG�u�4h�b���?!��	
V#��HJ�&��!LsDvH���a��C��u��o(�Zd��J����bh������K+�,��ךۊ��]�	V�]BN��C�|%�l�-�D�1)v1�����<"�D��>��r*�H�M�E��;�J�!��iU
<�X����B�5�|��i� #��Ou��L��9/v$d�u����_z���B��mW�%xU-��ճ���,�G�_��D�o������y��J�̙�p���N�_8N���L�Pj{X���*B��)�o�>4S�xE��$���g�Hi.5�<�	�Nj�5ٲ4.+��þ��Ɓ�NjG���Vʶa�'Ue	>�Mvy#ۻ������r�����n�xk��E%E"ye�BtY��m�eZUpkE�����ӭ�W��jՆ�ȓ��U�z�#����T����̃�C��4��)�����j�Rt쌉Čc�a�ZH������Y�ŵܰ�As�������P��I�xYGhIT#��vP�� �`-F�"�ti��2��}Ome��Sx4�5J����o8�J?�º=��.�kZ�0/-�Q�,Xd/�O�])|l��f�۬7�3�0����td�k���dE=�r���	�%%Y����Ҥ�W�Q��ès�(��~ ���8�����	�U+k ��Z	��_#qSWpD��*P3j����Q�r�IwƵ���n-���H���	��kQ��
����F�S�$�HJaLP兂��d��vh2d���\��� wl�������WN����r��qYC^��z�?�0��楧SƋA�Q%D�qϳ��x�$��;����
��g9���.�D��W���Ý��&�ҿr,�)���~�����H�g�XV$}����"���`�K2+!몁?�dx�S2TXiC!�TN$AEWC�Uj8���Y�����fTr���~�x��/�dR��]��U 2�p����f��ї�3$�N4��>J`�&���'	ӕ��ŏn�$*�$f��j!�Bvx0&m�+�};�2���]��WY�mKX�rߗw%��_%��rB���V��_�e��z?�^A����tމi�������Q�#Dh!*�Y�W��7>��+�049�(b)�k �AZ��E�ɻZF�	M[�Ȕ����U���?	M��\�4�E��e8P/�78�h�+C�:�uRs=;��Nl��B��Ѧ��+eIy�E#Q�:7X�dtL9!�h#e�#��m��)�V��_�W\v�lXŚ�fB��)	�)���	lMf�)3d����jM��c
qA�!�ف�[)������e'��C���q�/QU#�ՠ���x։t���]��(d`�	�l��E��=�[ �ᄪJ--�B����S��xv+!�.p�n@�7$�@�:�W5������KBd�x%��<���/v�*�-�E��J���f蔒�nQ/=tRCI��ҍ��  a �� o@�����[���Z��:g�}Μ�����y�R�f�˾�M#��ih���l4 NEhY�~ ��s�S�NYV���}�5�}����[	[P�_��A����t��^:D㇘��h�g[�?P� eG�f��3#�7����BǞ �q�&�[�p��ŉ`eK��3�l�?�7҃��V���E=RJ��0n��rYh�
��/�Ԣ1n��B��߫9eMOY���b�;bƺ�HxH��I�@��HpɅ$u��7��`����'c&�ߚ:��1�>��7�9�W��S�덑�:�8��[��օ��lΚ,~C�og�tj�WdC��Lb�#sĩ�`N��{�o�v,�Ѵ��'�+aw���x����&R�g�$A�7��Y�2�^rG����A�>$��[��\2tp� ��(aA�W��V����̧x��"��)߭���mȜ�=��LĆ:m�L�/]��+Go6r8�=q�l���G(�����F
B�+sޏ|��d�z�����W�UM���&���`���J6eӼY���ZN���X�_���&����.�sN�]lXF�9~�������_��F�.��̩�p?aN;-R!��v�rSxm��1�⩽��BI����w�6r�B�*��[�������1����$`�F�7l���4�v�ܳ)A�3���>�G�ꩱ�NR��k?\�eY�3)��F+:�뢚�>��Aސb�:���Gc�U��l�V��'��Vx��1| ���v����`����]`��,>�������ȩa��!B%��(.!��?��%��-�s�vbN��͛$(yJA��0sX�so^,���h�A��Ќ�S2|�c,fW��ߐ�w'�#J4[���ۤ+�n]��(�4[��Ol���Q�g*�l���O���FӖ3�)m��B�lNJ�'��X��[�<�9E)��H�c����4��p�Ԡ��_�is�T
��(�T��|��#)�֬7{�]�Q~E|�'g�rl�`� �8%_�O�����ipp]F���v^lF�|W�����"|n@�u~��M���y�ޝ��%8J��ѻ��z�w�c�㮦�e8�(4�������\�e���ZM���)�����:#%�4��/�䤇��Q�T�{��X���������3o����Js�+�G[�g�AcM�)�2n8|���]��Ds����u�}j�aX��%>Eȭ$�ϦCG*�s�~x�dsO�ҿJ�u�,�ʠ#ۡ��lb����d�*Z���������:�ȝA�=�ԙgR��$�9pm_��R�zi!iq���i���2��Z�:��&�wBg������/��t��)D;���'ސ�N�Z$�eI�p�4��7lV�����Op���8�C'P|�%������q�Tq�'}Gfk��� �j�0�c@��{�{�0h\��o.���2!����+��EMٕ�`��;B;\����?�U�i�dg�u��y��9��"F��G�Pk�[%'`;��=���H%�o��_ά����e��3��g��37Cۋdq(ϝX�eľ�ȕ��?m����1=�P�"'T�k�="�� x���^��8a��o^�1�k�i����B���Tu8�� N�C|���U1ٓh�Gϳ�|��̃\E�aN���<k}#�p&���*oϫ>>��ОѺ�1���43y�6R3y	����R	��&�o0��Oa��J���L��RU�V?�n�&q�\1ݻ$F�rgB�m7�*��` �N)�&H�ɸ�/B�/t[QZ��˩�+^6� {�~F))�Rit���8�����1�C�]"5��x]�;����#`��8d� ;@�����G\`��[��e����۶�8~ j>�t�`V�0�ٴ���;�k{��<W���%�\��tDڹn��M�}Crȓ�e]6��EHx;�ױ����w�	e'"�z��Y�8���O�$�ML�B���;��;�}2���p��AՏ�r�eJ�t���uA��C�c��9�/�Vy�J����<��+E@���B5V�Uus�Y���Cia?�cmc����i���)e��O1��&�m^�SBh�<U�6dyC�c�Xg�g-ەH����?UY�8x� �c4���i�ّ��u��(fB�L�ܹ^4�z9�[�f�:�_j���p�V��$a���n��A��U��?i�ei����r�%S�����^%>Ƃ*�o��X�b" �qZ��?�Nf-�D~AV�o4<7i�7��q945\[Q2<��5��}��m�ؘ9 o����2<cNUUB{��l5�Y�X/��E"�P� ��ޠmYҐ8�"���j�cb�c,��uj���?�@�<AÒg�b9n�m��f��ײ*´��oΈ�[q{����k�U=��M����3Eq��,�F��\slQ�� ^@�k�L�k�7O��4У�Ώ��̓��ޠJ�ӂ�2S�.���rd�|�֖�a��?�����RM�[��H[6������R}��Jrh�KҘɊ��=��E��c�_�`�/MjQev��X;e�o��X7���]ZK=���xG��H
1b�-�t&Ec&�-晖�g�����}�x�ދ�.�&"�9���S�s��r�:���J4ʣ��	��/��F�J�p�\nH/^����>��N���+Uu��e�à�Ԥ6��Fs�s��t��4g^*|����:0��NgB��2_�}F ��K��%�#�U��N����8�FKR����U��f��+���J���O����;��6=����T��_��]2�GI�aGU�j���kVK�"����N������&
߿;ֽ�w�b�kGn.�9�"�����>�o�<E��&��Ey��:�lwH�@:�e͗
�Z�����Et`z7vڻ������b1��s�U��g�R�{����A�d�����T�M�׮=]���9{�a�6ø�n)rK}�4'�[u���t�"O��0,;�0�Tt�ŵUf�*ig��3xi�����D,��˪��8�0�P��?��_qwZ����>Ұh���eo�O�-w��i��  ��"���G�u��:����	*="�c��DA*`�Sָ��O�l��}�ڡk�/��M��Z�u(k��7 E�nܸ�2=��=��%Y�,�����'���L����_Ȣ� ���9�4���&f};�eYx�sK�e3�y���S�V�|�yX�aDbZ,W�&����f���~Н��i�Sz����oBC�_eD�R��.��;A  �1j�<�KnS��E��l��տ-�.~�H�TBK�G�Ϟ�	
��ܳ&~��x�G�?�������]��r�W�ò�����F�v)�
� �1u�Qi6v�T�&���>�ګ���V��o@�vD�+J\���5��������������<L�"Ů�+� �d83QM	yV΢�k?<������)�����˯�1��ͰAyj@��r����v�Hĉ�⭚Yx^5Ez�1����l+Y{�s����Ů���*����#PA-px�:S�5�g�?,
������U�r�KKEv�j�g�}�;����Ld=µM���e�d�3���&�M�����`7�7���Q��S�]�gb�_�����ޟ`���C���L�ט��Ϙ��J��Y�!̢4L���7,�K��5:�㟛��.�WD�3��T_)�?x��i8��Y�C��ԯNIL�������%����^A���=�e,\�>��v\m�cPx���Tq�wϝG���Ӻa"����u;��J��x��V�h��n.v8\O>�J]
����̌Ie&�wg�kV�D �U�NR����N2^j���G�5r2�'��E�ZM;���\�m�ZD�Zc�������{"�_��~��'U�����n�e] Y�+d~��V�����E�7���nS�ʜG̢X���s�ͬ*�j�^
D�A�$���������̏���Qփ���}�){�Y��N���Ε�v��@��0���4g���v��}���Z��(q1t��"�E�'��Zӣ�\�HZS�G\�B���n��Q����<��}h�PS)f�^��p�b�dgR���nS�"ID����s�0�Z���g�;�#�9��̼/c��*�v�M�e'�x�U�jǚE���3�O?t�@-3a��KY�M��l}[�7g
�����?U<�sI*��%��@���O v���ݤ� ��Y�d�Dc���sB��_b����?�K�"���6ƍ4���e#��P�ě��Z8�b�1%|+���%�`�@�:��.#���1F�1־Wp�M�4�x%%�1���M�;�SǴ>�XlS߲���x��q���[b�4�;rN!7?�J�]P"�M�_�X����?݇k���l�Ao��JK�"?P׼�����I`\�7�Q�7�{b0h[�4$��U�6MzQ��c�d�>�a�$�X��2�����l����A�N�,�	�]n��Ю0����j6v��P�a��)A���Y����I��1\T�EUj:��mZ�-	Ud�=a~Tq�̽Sԗ�Q��Rx�U��1�upv����MA���lB(���G3FT�#n��W�""Ù;�Pf���q��v�#Z���s?'b���9�|7�ȉ��vJaY ��y���S�u)�\����0��B��p�,��}.��&/��lV�̽"z>�i����̛�%�aֆ�����w�i�O1T����|]%��
PL`\�t��m!-�L�L��M��L#�bu�;��S��W(i�y��:_�Ŏ����@F%��e�<U]����"��LtF:�5���iyL䴕��{}�*'���ި=ך0Ň���IrBP����u��^��0w����W�I�>9�������Y1F�cTM�Q(vJ�/O�f�����3�W�=ѥ�6樉��s���N�2������X���A�Re���[g2���>��}�Qb�4x��[��$�4�C�[&�2��I5m�~?ƾ�s��;�/xA�	?���?����s� �i��	)8(8[�oY��F*d���=�&8S�<��0E]j0�)�E�uC��4����x|���4�+�`�n��A����Rg~�>�c,\8�	g�UI���?�j��>�<a~:Ҋn)�I���E�o�?ܯ{�-��Y)�1�4��t}���ƌ#�*���_ FF��R��v���^"��sܴ�Lޚ�(qK\&�W�u���X����^�C�	���RFS�6w��"�pzYN��7��ŊDqXgvS�B)K-�bf���(ӽF(C̈" ɑ#w��j��V�Z�B��!�<c#��x�+n}�^���$>?��Y�m���N� D*uW��\�����ri\ۼۀ,(ҧ@�Fk�p�)(�s��V��p��i�����fҰm._��&|�^��w'}��F�x�4�ANA�,��Q�3Ԇ�h2�������b��'!L��m���rRM�~��)�y5 :P	�vq;�a��a&/�N���!��ئP6��D���_ūvPq�wy�ލ� N6�ᦒ��I8���dx�ӣ����!ɦbESi�g�+M�!�庂� x��1h�N	���R\+��F�������&z��&�q1�U<&q�XY�7k&zM4ֆg�+jb��#mkl W��x2%����P�.���l�����DC>��~�:" G���[ku ��n�����d�MÑ�/D@���Y犘uoѹ�6�`��i��H�k�94���p��D�� �٠-KR�
�F_�gb�FBI ZpO��������PɋS�%�{���� �!��^
/t�	"_��O	�\x��E�n�����m�|��R�zս��#ӯ��>@�_"b���ު�z�`��j�64o�Fh�����h��OO{�<jZ*'���iu;�ɼJ"G�
o�N�ɀN���	�}��c=Y�O����	V��E۝x4����yÓ�[�n�8B�`��������y�:�A�!p}��?(.��7�����އu
����m�R�"lǔ��4�d`LWً��}�qT�(>���,2��L����R�K5ՠ�A�
\ҿ@Z�H��BI��2$<k�����DNl�4� �򀢙�?�6vUQ�\��WY�D����?�@�����T	�Rx��X�����F��t���������yk�W�����Dcm�MF�fZdE��bI����op�d���u�f��a��{+l�*�C�3z
�f�J��tc]�>c�oZ�.(�
�;�E��PA�J�L��繟�э(y`��-K*1���`�(��ʨ�%!xd�mA���I��`*�Á��+�^큏�P�(_��
�g�޹����E~�6�;fo�����b��]i�a�A܀�&���Ȼ9S���_��Ӑi[��ɷ�ְe1XSg�r|�?�tNx�f�m����KUIG6�Q[�9�G���k�s,NN�)����E�o�/(.����C���%�Dʩ./6��?zL��|�'��.d�.Bm���l�z'�Z��*)�TV��L�#�p�U�6gmt�¿Е��%jb���q���>��J/Ufn#�^n�t-E���^�d$%�f�	���Z<Dg�f]�*���$J���,�+�>�=��1����Y�{���F9>���o9q)��R�~?��x)UW��~��I�R��	��_.4L���&n$���R,DÛ�j�����z��Ԝ#�iLf��w���q:
���R��i�a
���#Æ��������[�j
x����%����:��nG�a�7��3��4���i%ξXFҲ��@⭇;�?3�c]�|�鐔�+�Ջm���.�{#�,W�]�'��ǉU�هM��z��_e���}۴�L���f��)�-i9c��m�u��\��蜽&y/|���<������a�C�ڢ�����R:�<�*�q�zy_�!��\<O��;�������I���g��ȯ��ߣ#�I��=��H6�n���ӳ"��p��]4���p�Y��@��cd��Hwe^�?��o����V��ihC@��:.�$t�Y�o�?
l�/[K��w��?m��Cl5᳕ά�k����B��0fB�S���������A�}ͯEyhСC���u{I`����3.��Ģ1=d�_䠠�Z�ƹ�/X������H=l�=�ģ���J�2P����9DI�����0��R�فvi!�S�oF�.NI��N2s3�K�Q�p�B���fN��Κp��!�v�z�,k'�\�O�Al�+s�[1l��V�_��a�Q� կ�����n�cm{�	u)Q�H'.���H���@VHl��F�5�����;"��[y����Y�CIo�5�Z�ҍMp�����6U�f �����g:� 4����E��i�y�5��P�3�)����3��
�0���ǮhtEM�\���c��n�.7��;�T�`��@���_�(����l@��ʂ{��m+H`���/q�]ٺZIa�Y /ܟ�%�� �S0��[2����R|B{&?�^��^��VR�����$��Qt1_�]f�����fUp��ԝ���H�"�%T�)# �?F��:�7�W�Z����F+�i�H��Z6Δ͍����V�Ŭ�8��
/�sH:9.��h|-YZa:!|�\dIJ��K?�hP���*���"�������R�M?��ś�VѦ	�p�^itm�v�&T?̙fap8�CBW����*3B�������l�q� m3��1n�bb��k;�F�XW2ː�1���}q��ޚdFw'9�Ü��*�R������F��UtS���.���eD%a씘)F!�р�+�+��eb��D���Wz�]��y��o�q��E�V�W���am����﹐�_�/�o G�3�nP��'�ε~N��t�<C�Ћ�S{Y�sk�Q.|P�E��F�$\`����^�G7]aԮ'?W�}��dd�̇�1�[�#����$���æW~�w;r�����T�Ұ��\0?F�-kJ��I[Y����&�l�E$��OCE^��3������o�Ͼ��)< �m�_)�J���*s�4U�!{��H&ϱ�7)�Π�6�v=Y$�m�7��&>Y'���e�l?<#�@.�,@�z�]�D@�?�iI<Q��E�1��&^�R{�/4���.��|�<�R^5��))�2�j0��.o8g�>2�j�2���A�l%�K`��y�w)�j�q��T�q���aq)6�ǅ��Y�����d�cS�I��oF��O���A�
�Vut8[�t�Mw2�z��g ZQZ��ݐ���s�0D�+Vs�#�G���7��ݔ�P~�V{	�uta�`|�U�1n��Gf��0O�f�dQ��&�ö�.ɫf7��w�2*\��ns�|+C!�<�����&]zB�Hvɞ�'D�EW���\$�)%mg����� >œ�Ei�o�_��4S����3���_�_��O��;r;��@�ЩN�K;pR���0������L����Ǟ<R��"`rs}w;g���B�Z�82N����%�^L����撎d����X����Udy�Gu�S)E��)�
4�.�?n���VN�;��5H�B�p$y��	�J	!FŸŗ��7`�0���	ϭ�=+w�=���O��������.[d!�?�6���'1�p��=����
urhd�h�L������x��l�s7.�em-��e���4ʰK�Ne�}O�r@�
Oٜ^P�+D���P�l�G��gH;8�b�|��@$�Q��ta��Y˥+
&>P�y��]J/�O���n��d�٨J��C�V|�`�F��k���Sp������`�f�t,̅(����kbf�CA��Fr>o�{rР8iP���V77h�]�W9$ �j^KL�~����~G��e��dr����*;b�锯6���^�3R~DE{DE(=���A����D*lDCw����O���'\�g�x%�L���#�����'0��f�<�ߐ;c-����݀.�j1�]WХM��selö%��� �O�.��;��+�;�p��Օ,�>��P��:�[����¥��/k�&���>��"��ښ����X��.�ȗ���OG�G>�P��;s9i�
r����V��%���`�V-[@���.K���m�
��u��Bi�)^Ƚ�̫d�ô�W�(������'#�ҏpR��{%b���%�i�X�W��p��bd#@�-��D+�0����2����O��G:�g_�^��Aǫ�?g�6� =b�H��'Z�� �Af$�H4�\Q�Z��
���(�R���7g��2��G#?�]�68ݼ;i�d��%��USJ�j����3�<�B���,kO�ފ`�93�fq,�L=�n*P}�8G�sYkc�l�-C�x��>�*W�G]�H���`�ָ4o����\�$�"L��@]���K��(���� \�Ȥ��R:g����1��#M�Q�f��9�۱����N��*��ݖ+�q�Z�'��B�(��fx���y��Z�Q�1粙�%{�����R;��D;6�F��H�l$��>�����i̒Fj�K��d0<�I˫� ���L1�eVJ���㈫�wn�H2�T���;˘*��k�p#ijIK)z\��'7y��;Ͼ~�~DS8��Y��g �Sս������oR�#~7/��n�K8�sOO5�ڭ5���,��lN�b�e6���vw�L;��<�bt*�E�>N�w�f�JؐF�1V!W{F
��'=�^8��s����2�hCkM�t��^�g�"a9��z0��_4ć.�á1��(b)�"�������t�
37���ٰ�����ɻ?�w���Ҥ&y�9#���+(J`X�RVn7h�dX�LI�{�a�s��L��J�����[L(���!9@J;�:�H�ek�N6��z3������w�ma>Gң�A���]�n ��p%gÅdس�H�>ʦ�OA�Vd|2����W�t6�����d��!�?S|׹�b��ޒe1��T�k�V��9=2y���v:�� ���Z� ���D���d��ؕ�o��W��G ÷K�(ؓyQ�wG�i˔�����4v�)���P�p�0{���h(��j�����B�C��&����5 �OϚ��VX���ȃ����n�T�����%xm��S;Ե�7}s#�o� ��x�??'<��v�~��KUuG62Q[�7rF������hDΗR-���f�wv>��ž�VFI�P�;��^�F�C�����؎)��󢒩N�RF��]�����o3�����#٩��6t� �^�|�zԞpM�^ʳ+��Q��x�2��w-0,��3x��Ak������ ��y��{��k�W���<�$�]��U�kp�䱒��u�ю�!�N��N�qTos�S)�K|��y��f �m�%��ߋ��ZL��I�Q�Y��p�q!��
6���=J�U2��+����K���|d|�[}3W6�H
�K�C�m3��RlX���H�����w�2QuB<e��F0��n��נ�=�4i��Q�VO��P]�镹�"�㍞����l�s�w �8��	���%׮�䉛v'{PLXb�mR�u������Ga;q��
��_��Yfx'��)�uA�	u��F&$��H�fW������6����w��4�Z��d� ����Q�奱��l"��#��"}��zz���~��L������٧��`��BK;r�Ԟu5���J˲������nӳ|s'�����*��Jv'�69�[�U�X~��Ͽ����x�6Gsv�N����F�ף�:ɢ֨뉣'D9)Jv�hXP�HN�_n��n��A�`t��Ӷt'g9���0������F�EY+�1��ˋ7�x�S'[J�a=��.Q�s�4_�˦��}?ϱ��f^��+���v	����+O�̥ؔ�g��b�(6�����}-��ux��`h|՗���y�a VV�xg�Q"e��A��n������~{�2��>����? �~Q�5z�I��`�~�L��@��d=|r��d��`���W�5�޾O�6���q�O��a������kD�����_L�|ѓ�}_���I����:�"|$zgC�u��1V�_&�=T$��� [�k^���|��^���Z���t��Ǌ�����D�,��$��� ��a؅3(\E�/
T���4<�w����4z���zJ�[ �o��]ޑ��s�����I����[���ȓ��}����ϙ�Q�Nx�u=�B�2Q3���_�P&�d����!��1���G'F��2��^����$�<X�Z�&0f�����ߟ*wM؟��P���*��r�~	�(r��k����_�>Ə�"�ޞ�^m�������G���ST�'b��i���Q��A.�Z,�h{m�����N#����o���vZ�6���F	��)��g�X�O
B�bt�h�L��ʏ��6K��
��I���/��#��]�&�I/�oVd����ؿ��B���v�K�����ZJav���'�~�3�d���0^õ����O�G���>�^$�h�.�q��mq����Y��ٲ��l�[�ӷ��!w��t��fu�򖧐/ϙ�~`�M|9�I�s�L���nj���҈e믯c�I&��r����ǈn��_�`�,o�>G�����Y�lU�aѾ��Lfd��4_9�ZY��1n��,��+��Ӆ��w�92�v8]K����ǥ��%Ӈ���J���*-JF>�)n���=OI��U��wz��#��,_}'t��s|���R!�k<��+�)���_�q��ړd�oH�O�
����u1�T��gUL�\X���tj��2y�����w<Xկ>lK��u0��H�"s�O�A�l��.j��a�Q�V���̰�k�=h��;۪�z���޻qS5��Q����j������''�!O��!)���Q>Ĝ$ f��Q��k��|'��-�w��@���7��|�zk�A익���������G��E���$��y�-�Ϲ�"|=�����V�G���;��z��>V�e�x������+�xV��e��y�E�
Q�Hm�ň��X4�ӬY�;oW��U��.�QE~gŗ��?ocDBnR�{*o���ό���$k���%��L��o��7���nō��R\y"�󕝒ރJ���U!uG=��c(�"�S9��P���g�wL���J��@E��aF���>ʏ�r�I�p���r��kd.8ٖ�k���/�"<J�6\]��{0m��"F�9�+܊ՙ��Z�p��-̪�:n��_�	JTa��])Y-O��O*ħ�)�{Iw<�ao[�k�x�#������9���SFs�f\Ot���l��,�	�f���l�W��&Z%s5i�k��ɊOՐ��M�&E.h�X>IQ�9Q�I;4���0�w�d�_�z�����t%��9KgG������(�"PJ.-6�t�%<3kۡ�m��/�iK-E���!��g}�O�	�����9��h�T���	<�;i{��}%���ޡp^�V#k#·�hsR�Ʊ��9��=�)�3�9-�X�h
+���=��B�g���n�x��n.��px������L`�����3��*���>�G���8��uQ����M4�V����u��yl��Ν|�0�sdB� �����W����e�vHג������|�t���T[_��A�x��z"�$I�g�شY�d˴2s7 cwG��S��1c��a9�3���c/�Fv��kʄn�}J����0+-��i�{�x����C�LU�-����"�2��H,�+ND��3�
~'��l�&O!O#%�x���g]�|����e�t��;�Rx��Z˅��[�y��f[��*إ��d�/Z�.7Z4 8"��$cZ�r2�v]R�M̓>l"g��_�}�z3Fdک���/s����]<��~J��\��e�RQ9����D��sdTD^Y�*�z���h�[�x���v�u�uYWf��X� W�	��=Fzg!�NF�É�a)�ue�U�t�o!�P��i��Uh�e�ڗ�8��c87�8O4�#~��)�ؼo a���J�5���U�wُ�����G���
L��JY�l2����bSN���
!N��r���r��!q�5&k���c��x��X}��X��^�
d�Go4Ky��(*�����.����v���$k'�o
�t|)�z�������Ǐ�QqW��`�B�,�%	�S�q�-չ��~7ŷPY���"�!����/X��Z�#9����v�Uz�֜2�B�9�E=��o��^oy��m�g�U��U#��+/~ҥ?��'9l�:�ɰv����9��u�A�(�l�pя��nġ^�U������:��ĸl~�'Ψ���D:(��g��Ncj�Z-уdX%�9c1�MĨM�B$���z��
�LU�� n����7�Ƀ�麺�X�K��jf�#�`��۴8�~�_�o���ɣ ����;�T�#KSoY+�X\mTI'殽xSM�M��윆�̂�\b���L^^��ZtRW�QY( �����b���e���)}�T��*�)J�V�0���Z�J����|%�W�q��a�����E��ǃ��I*���,>^���7=�J���>X��/9|M*>�h��({Qy?G
����^m�Q����^�>�`^�U�kD:�up|�W_l���Р	 K�;�����=g0��Uu��ݑ0�U���t��J�nF��xI}�d��y(��d$�`��]���2�{�9�|b�u͉��|g�H��b�b[�+qF�~SrQ��OEo�����?gwet�&_���>����Q�oȶ�O%��4}��_Z�9Ɗ|Ҿ;va ��H۝�&Xy���{*��,�c,�!��ɡ�[���#6���۷�կ��
���w�D��"�iC���-��ѝ�"��ⷷ(A9�H��� ��i�s�	���ی�KJ���
�?ޤ���E"rU�=­q�R�qK���m�������g���T9ة\BR�Q�z/�����އ�vW�M� ׉����]F�m
��K)5�6�ʶ���-s�T�pqEZ=�Z��%�IQ㛫� ͽ�*$ޫ�`�� Dd�&�ۊ�<�q��k�H����0��9+�9Ww�{H��x|�Gw�	��!�VB�{b����,t���NV��2b>�쬸�F�b�ea:u5��)P=�Q|��m�G
]���=���X�#<�KmK�����hاQ,�@�X��<�x�����*}\��������ڥ���l��d�@���a?��*<UB)�Ϭ�񃟼)j��ӗ$�#x�f���X�;�m��X�E�2>`�֢�������-��e�~�����R��/�ט�6�D:k��)YT�M�Ss޲�6kG��g��Z��؈YY"���:����+�X�q�G�Wae���E��3����n5TՇ���/x�0�ÕM��AD�!�h�u@�M�Ǎ��ƨ�����B�@���@�Nh1�����y�o��3��¬9����j�^��Y:���(��18oc.;�Z�TTl�ʕ�v�d�1��]A�*X}M�7r��s�.�A��@ǋ���+�v'_���z@��A�dr����睖��@d_B��À�7Yk�ֈ�cϚঀ6z�&O�K�������G��t�����3cJ9QW��騤:��r�-�����8������q��~���#��Z���m~����Z��l�asI�O�~�B/ELZ���f���f&roj^=���&���_����]��������� /;��,��c������D��%����Vt,ѫ#4l��)W^��:�Q��hDb7����4�gej?z�^[-��d����`Z�7n��s���� 明OEQWh�K.ͤ�Pz�f��_<~�e��&�=��MTӼ:���`H�9�
4��s~��KT�0�y�L�k�����lĽӑ���p�Ё�ϕ�x�M�T�{�c��E�)�üm8څ�ǟ��l�=�fEt�^b��/R��!.N��o�=�SUZ�%��إ6`�n&��[G۝ŋ���ɴ��}��['k��T�����%���H�Wȹ�w7�$6�v0s�Gv�%F�q	:ʎ�$�o����tw�FF45y7谮�\��t��!/��T����Zi��W��I��A�R���x"w-n�4�4
�����,��VsiK>2���M�Q���8rC����ݸ���T�Ƚt���!xZN��{�dc���gyz_%�iM�jU
�(/�iut����]p��W����4�D��XW[N�wb:��ks��e}�m�\��}`��~c���x�63��^8�)T�z��x(%9C �M������E�8��Rw/b$F�-EM[^O��a&P1���!|�5D3_w���[#n��H���������>��Gx~���08��C�`�j������B�-B�B�!%���I�9��fgl��E�8i#�\y��;�U������n�P��TX��ճ�u��� �>䷵(���y:��yq�u����|{�ŽY�����oĲ�*Ի����|��i�GU��zt!�ߥ�c�{�
#��O��w�Y�q���w���:�aP��� w?x�/q:M�|7��W9/��dV��)v��<�(j[�|���\�ToS���i7#s�<����0���;��	���c��a���w�3�T�c7j^�4O�I�韠���9�~ۧy��u�ؑ��D.]6����[s�6���{���ӛ�u������f�n-
:GQi��<R�E6����>��ɲ'�M�'P��Vw�.�ۦ�����cތ
]s�xP�>ۉ���B�P�����;Bl�R�{*�矊�L�HSI���됋�f��u�3تzq�3l�����ۋ���Vj��T>Xd���C	�R%*����MMb�z?N�7����,����W&dZ��`=nvWJ����n��Z#�(r�&{Z�x<f5��2jW���s�w�=�z��vӬ��`����+��7!���o;�Om\F�T 7���XR�e�4<�P�x��;�/1w<Hs�^���R]CV��2?ʨ�a�Ŋ+SD��8����>�G~��}��9E�����6u���LۢwFA���8�x2�gO1
;��
�!`/�w�5�L�3�-�KvD,ay���>5t��ʽ|]Ј���ހ`x�*�6������x�5^׋�w�k\-]�C���j�ʇ'��U�x_C-Т\���p��l�%���$�Q�����'Y\�5���x	t��W��[�!����553�_�~
��n�#�"�J��g�l����KynV�<l�v(*���P��C��Ƀ��Ń��؟�)�Tߝ�0�q� �܈ �['��	f�:ڤ�=���u�����H�BE
3��h%c0O~H�N�\���M%����p\N�����)�*R�<��*IԖ�W�A�ۺ������՗���˽~˛*�i�haps˄�*Y<��Ϟ�p�~�������9�y���Lna���g?|��5`0k�d�Ҍ��?9��h59[MZ[�>_�F��ϡ��v5q�BU%;���"��)G<�M����njD}�m؞��+�vK�{��f1�ʊ�#E�g/[Z=�v��\��n�\J0y��xV���iEP��|���n|a\�H�e��(��A%�B�p?�gOJ_���f�M	��B���mٚ�"�wڻ��>B6�m��=�q�ّ��KӚ�����4�hF�V&=�Mx���b$�b�8�5�M���'2-d92}�e*� Td���px�U|������YF����J�Q�3�JN�i�V0��H���������f�c����KXgSE�y.�8F�"FH{��hO�����$���߬����"���S��i������J�B���|��!��<Wg��1K+� ��"�PM��FH�*�vs� ����t*�r��J�̶�CBlwoF�nئ�"V�K�R�������|`_X��R[���Z�\p͗b~i�j��%��G$Py�U��!� T �{M�Y.��֑��h����'�.j��W�C:F5i/)���_R#�ѭ+��_Y]|�A���%{�<�v�^p#���O�P"�i�cp�5��K�!3ƒT�`j�q~-FN�,��a��a�ژͷ��:�?��y�� ���?�f��TM�6[g��5��^���Q7��	�XI@�1�B������;ӻUmx>5a.b����b�f���?�w˨���m�qwwwwwwww'��@pw��Npi��-x�{B� A��侟�]�Y3g���}����]�w]�޻�	{Q��ͳ�<wmù�!�/�}�W�	A4���l艿 �x����B=��%������-G���m�C�֚�鎯|�P؀	a9z�$y�>�,ҡ5��`,�;��y,���>�wM��n�
�0v�7��E�[�M��d�a����.4j�����d�07H2[��`�����A���m�ݞ�if�Y�z������g 2c����7A{�.�JR��p��R�S��f�Al���F�+��� n%�9�XׇϷ-��k7��|-��� �v7�n�xI�VJ��3��l��o<�<�ib���UW��)��tp�A���afۭ����U�i׸j�e��c|O��Q0Oh��xH�/˺!hf�a}���8�/ÈI��$l~瀅f�SjF�Y� �)�S�2���?�@����DBN���%�(��=��-�
��/��q�-�*�  ���
*�����BN���ǎ�xc�}��@��
� �'��Z�z����-X�9b����B�+v��>��A�塥7U�<����л�����k��Rp����.�9���B�˽}k�Ay7{7
������B���M�[-t~�!��~��h5��JU��hv�k_c�����"�v��V�Fv/�V>��å�TF�V���X�JW��ow��S�s
�9m������}���ˈ���t��p$p��.�m�7�Ã��P���p:_!��˽�M䭤�S�8�9��"�7� ^�Sr����m�k4�5�Y��\ٙ��W�	��:�3�� G���:��W�.�ҵ`?鿡p"%��)`+�i��¤���DF���W0� �ȑR�ivw�Ex7���cY�J��W�,�㵭�I
��|��ԱSI̝���Co,��j���'��wH<zG���XW�ƞ���|���Jɒ��������"���A��J�C�Թ����x6P��O�2��F�_��(���py�Q��s�������U�.�Rb�>`c���ӟ��_Z[�Z;���wR��JS�~764��6B��D�A�qE4RR��&�w�P�WO���)$[¦Ow��>�wЖ�6�����4��G^�ܘ��ؙ�Y��N�k����DM"����'�*�����әJȃ!�d̈́����L��h&50<�P�x�f�)A��w�@Y��(�okiK�3�boS��/����b�&�\E���Vc���\�U�4IQ�i�}|癆�;���%)�R�/�@����Zv���U���t�S��v��o�~V�Ρ?��A�����֟x��`l���� ��.��|�����P��� �$����Ɵ��'��KSэ㵲�5��^!5��d���ׅ8(N��~u��Y%��u�)@MAx�`���45�CǤgVQD=�ZCc�^�=��_}��X�+��V�π;S��@�su�v	[aݰA��z��LNi�FZ�44^>�����c��(��1J�!�˟ۏOF5���Z��(��T�0���N��h���k~q�E��l�s9��a>�T+�`%5.p�y)�;���7���J�nR�a[�r�ՌV�
K?��԰���Bva�1�����xe�A<�=$A�|�b8%<�,��^օ�]�J�߬�E�@�(C9Ml�`2�øa�L���C���4�9�Ee�!9�I�l�f|��)H��H�UF�M�5���q$9n� i=���\þ�����-<0N/ӓ�5X7�����<�� k� #q�Z��v����[~hr�m�-��*���H�6�+O�+���b���m����1<&�s�W*��ۓ�(B(X��Ԓ��o��=��2���=4r�Ĥ��?�4�}D�|Gp�!}�3�w�&�o�͟X� P�2��6��-�&�8dbĺ��@��[h�Q��F���2&�U���� �斂v�}	�$K��?p��ǘ�b��;�lyB���^����M׮<@sW<��z�����D��ۼ#�~���J&q�����1	�'��:+)*'���eu�H�a�w:�����O���zb��9L'��s5˙{�ZG�&�U����s0̹=��X�t��6+�Kd���e�*|�済�$�������z�
;��U��-��zwIA<�iĝ���,�t����P�m;[��S��5�$h���:�A%X|�+���M�K˨8n�0�������aX1���,��|md�O���	�G�<��OX]��g{-�h�Y�D��V�1����%p�Yh�����������WP�'%���_?OM�* ��wvM��М�����Q�T�<5P̈����m=���A֊Q1�-(]��}�61�^��+R{�F�onb ��ߨ�U����?��F�ݽ�9�q�C��Q��$<t���Ð���Q�����$1�Z䶶���yɯN(����qr�(��	H�h?�)2��lX��v���k/���
<˺&�N<kq���s�h�ᎱH�t	{��,��+9�N����Ȧa�BR��˒\9>\��NX�mA�A$�ni�bXd<r�Ӏ�U���3�
lk�4��{!��,��Q�&������ƀ��D�.o壯��y��a�V%� �g�vY��?H�t9�#W���9ϊʚ���9����&]��Fk�b�D�dM\I*�G�O�Q����c1P�)#�A㹵K�V���v�D��"f���'�Fz*{<�K���M4���6��Kv��rc��+����P74������f�C�z��i��9$�N���v?�K�C���]"�5��B���6�!���G�-����zO��M�e~�R!�57)(���~x#���/�F���ɦ���3A��v��L0�z������@8`S�RM�ß,)������oz�ɁV�HaF �,�ǍVQ��P�)}��Zy�􋏗ΰ��ȎBJzI��͑1������w2bٗ$u��hemAHi:*Å|��6j�	���B��K����c�h�k�����t_;}�(>o�8�ij��㬷;���/"�C#D�{Y���50�;)�/՞���1��Q�J��l�[ie�m�OZ�/����Qs��)H�
`�j�g�zs�MAE*������3Ҏ����yv�!V�[�f�;���[\i&j/�or���<Xr29�G&p�A4�o��z ��	K���>ￅ����".�CY�k�#��^�I�%�\��y�O� ���Y��K}���!��������]<p�Ff��a���RW��W��l��E�CG_�SDj�]t�"F �ShgYarDtS�?[���R�,b�J���k�X��ߠ�]X�N�V[L�䂓m'�e�,a�����*�M�"�4k�(t�aڽ¦��L�����kbF�Z�>�����D�pɞ=`��SHx���s��l�`y�]�����z�����`&��(x�La���#/;f�׺wF�9�N�.���蚖�2�:�"��~ܬ��~�������/��l�UhkI�dɡ�u6��S4*��8�t�[�����j�iAz�ى �&�@�w1�!�^ ��߹s���^�f:�^-�8TWGS��O9��
~9��� 8{��P�eU[X��3��U���Ov���[ �K�%���]�H��{l��I̼�	�`"/�������I ^{�[vD�hɶ�p7Ͽ�R�I/��i\}8�S�'#��m���
�X+��YYS]��dPj!1�?�qk��Y��h���>�z6��$ԍ�<��]��C�k�$\���c�%��(���B\Ֆ�N��7���ձ^n~��3�4�k�G)��i��q�o�	Y�~TS�f�#
F�P��%f���«���\�5�}g2!��>�K�(�:>��]�J�Ƕ�
��������4TQ*P��#� 6�R`ׁ����G:�0_;tR*l��YE�d�+M9�	�K^�Ql�ˑ�=l��gY���os'�����վ�ȋ��J���
���'�L��l"G�m��XV��9��2bU�����#�\:]Z, #!Pr���AF�ir�O��gӫ���&�!���gevz��>~-��BAo�r��W�lafa��2�"t����aw:=���W�`�f�Z�N����Z�l-��%,(<|k���{��Z���]�3��MU���\�������M�󯗮e������������|n�t�ژ���`"<x��~Y\#E>%x#����#�:#����ܗ+���~�ң30�?�j�s��%~��9sH�qo��y�g@�
1CUS99|��S�
�RR��cT�!6o���@�♴�鐓���6�芾�S��aC��v'���S׻���(�"�$-�?��=��z��4�~����i��CNL��S�eR{!������3�{�x�π5�����7�/b��%!6Gȟ�0po%:�n1��X�m�3�?p���a�p�
���h�f�R�3�rroP|��\�����QM��)7%�i��d�B ���?X��Y��p"��E��3���Z}��,����h?�E��;�����:*U���/胝Z�U_nZO�3X����!��PW�	�{���ץ���|�Z.����_vT��\�����]tW:@
�x�ğ�9���n�����e�qﯯ�;;M�7��v}�j~�C�����H��:+���P�礸9+�|��d�8�~sv*%������+vJ�W���33C�l}5?��,�u��'}&x�֫��+:��� A��P?���91�d9���-.�������g@���SWLK �Ϫqe������6����p\۬��I����e�Ѹ��l��c�Oھ��?OZ�{� fC+7t��?�C�c�{��.�&_�%5F@��=�R�����k���P���ѣ�����ê� ��~�9�$�O՟>�axz��U��y'�)�"�e��ժK�QI�I̽.Z1��?_�|r�ap'�qg|���S����~q�%������v�st��62�e�^/��|7�pі��;�7R�Kx�
Ư;ݨ�0�Eo[��9� �9��1n�ƸT�b+�����h_K���6��=��46�0&Q�r[d��e��#A��C��9�M\7���[85�a�w�fe����uT�n(	f3�����[_`�����,\�y��R�=�g���̦���ۑ{@��pI�/�S�,Fy^	��ZFW�O��������m�,|�_�ѾP��M�h�@�������8�|Sc�s�ɒ��'���w�ML�B���1ϺܕŻ��j�O���N#=�;�0��z����d;C3�l]|ټ�T(�Ͽ!|`A�bޘ6����h��Lf+>3.>Re��z�;}ջ� �g #Zp�p|.��Q����|�����ȺGP=�,���F��!m(����8�oY�{]�Q���Q|�Cgr2���^C��w1�wi c�|�ep��O��6h)Rk3&N��uF�"�-Z�sG��!� G�Vg_������4�s���!~���sˇ|�O��Уg����>R��XN�B1�s�Kcru�,駭[:�w�pr���ˋ�D"�<a��Z�`����Ƌ|\[���K�.�?7��L\}"��*2΁�ѷ�x���>�GSnn�2/[y4�ҦG�ǃW)�:��b�2�����k�� �t�#��;�[F���Z�he������ȐQ5�4"F\v8R��Z�?���M�H�B]y�w�����i� q��6V�$q���?5������Ai�Ό�������"Z��e�=���Z8���IE���G�嘞�D��5��;"G��tP� ]OK�5��A1O�#�s����Fɷ��-#MM>C%g#�t��h=�H���o� ���b7lKF�|n�P���O��"Ia�,���@oJ��e�\�=Vς��^7|��59��00�b���~�I��޺3�!?fA�y�;��XЩ��ޢ����F����vm��>��?����W�AQ���as���k����'7^��姑��q~
U�*^M�����z�S��P�?�
�����~�{��!�B��V��Ň���ۭ� *  	����uQ��J�VH*�f�z�z&��dڰ�����9�X�ΎeB���:w�zPZ8��6�}��r3���]g�
Ӟ.�����3<��6��2�i��>�w#� �b���la���CKIW��7J�{_26��V�����ئe=چ˷�g�t���2��H�}7 ������S;�Fp���^�����oB���`ހ�Ԍ�k��+Ԍ9ui�I�dpyJ��%cL�x�{�b�_oЁ�+�qjDz敵�ڷ{n�[���6�i���l5�%s�y
��^��w6g %�ɰ
;?\@�E�W�Z�ti������<4b)���XV�����b+��K�]�z�.b1 ~Aԓv�*-/ru�F�T���}V�DI��y��pV���Ո^p|�g������� Flp����4}��ܘ;9���a3�2��I�2�i�zԍ�H��4��&M��̟�g�q�di��A��`d��|�d:֖gX�L�����f���Ę�|v��ً�Jɯ�����3���	6�^�����geRIo����(�\�S��l����bQ1� ��0&:H�q���y�i�q�K	X�%ܦ0c|�W�]n��)�����QH��+�ѕ��#"\�C�k�s�bYq[lɎ`Ŗ���n�PͿTS��O���/��8�r��A���?���I��f*ҹ�x��n$���Pw�S�v�h�e���	���i�i�[��&EY��e�w���¨5�����V %�b��:),�e��2yO�\ن}ȣx�W��3��%ý�NZ�'[ũg �g50m2��,�=��֢QT*�!W"2��(���ňo�������=a�G5}�����"8�\�����m���?E�p��Y9Gͻ5(Y�w:��C;�i�#�qċ�6ʞ�	U�R��j��O�	2�ݙU�BY9w��q��4�	�X������_#��*���_]��8	�6�o�IKh�.(��
H�H>��Z���)���cj�3�$��5�9܁�UMON,B����e,��v-_h� ���]~s�P�
�sC�I�Xfk��v��0���KV�����u��C�����/�8�{���E匮g��Tvg:���}#�@�HP"��9�sb��K��p>Ӊ[d�.�:a"EB�p�~��-����.�
uI�
���w)���D<U�
��E�k��UV�"�%ޯ�o�� �Bv}�|�9�H��ov/wopk��͈J�IXon�Rqݏ�U_"礪P�����a��k�rH]�}�(��+��_Xޕ`���;�hY&3�pӲ�t�.?V���Wǉ z��?85��8�GR�3�#ܙ��'S1��a9�8�Or麏��.�.q`�3{P_Kwe`��䈊�]�@�:�'G���@��|L@q������ ������� +��X�Zp��������1PN�p4��`�F�Ydw��P7\�C�K��B�D��6M����[�9�j������� rI�~��ʋ
��4�a�c�<�"Y[��/�Ϫ*f��!��'a�;�ػ��}�̈́�N�.���s	[������ۡ�!�Sr9���2M~I���Y�t���o�22X]��E�^��iB��	>�f%�}�"3��fb�`�};u�(�<�e���	0�У����F6�Ò7}:�����Q�r2f&`"ۜ={2������+�Ƭ�ic�7s�oϾ=�])މꆻp>�a����@E�������Z/l��-Ս��K�]�+�Y`�,.�ǴGR%�Y�R���A�>�6.c++�\��� .��F���f8Y�l~�`��P�Y^��g@1��uӘ��
jT]���٧�Cly��CՃ6Nm�0*üH8�z������*��E����`|r8%0�d���'����X/�uM��4�_D��L��q��0��g!Mמ�M�/J�ޓ���/���ؖ�p�i�k`A�'aUX�T���[C����
5}+
 �"S���HAY���Q%�((�^z�4\�h����T�O���	Nz��lGL�C���� ��6���`�U��fS�Ş�I���j�g�Z"0]�I�*0��0+{�4`�H���}Y�)UM��;���{u{�㽎������/V{������,0�	����f��,�Z��g����5���`S���Z�h��G6��[_��-��%�3�P����!tPk=�|Z�y$��,��Py�ik��mQ��Yˏ_�X��X�an�rf��X��%z��5���K��Z�+�e���w�����bzH����/�����T/�h�K��O%.1��~��[�6�t�lF�Ԙ�s뙲^xDx�Ba����cG�m�N6��f���$�NJR�H�3�|4�h��o�/T�t�2�Ŭu_~e:'�c-�yV��ʊ�r�e�Ǌ���[�4;�X�ѯ.h����e�l�vS��2<2s��ds2����p�ү)K��i|�:F��U^��!%֌'����7��n���W��G�� �a�~���3��P�@��ߩTLt�.��*�/\�p�X���dqA/���Ax��lе�R�A��ۘNmL�.u��Gde�
��,]8vr��o��:�x
V��u���d��h�ٷYsAHI5��W E��8��ۘ(�T>���oMDxb�z�r�G�5���KD��m��l�W7Y�l���!enge[��B�{�������.&�S��~3��j�T��V[˼�]�o^�I0%t�'�7oV�M��n����j��$��$���1Du&[Ʀܲq����$��2��1���B�^{���!�C�����D$�x_�y	I�0��]�:i� '��(�_K,Pfy���WÀ�����Bi�����8!�ᓡ����uz���]�~���h쐿����Xί�Z�0�M���J!u���/�@c��#�!�nƙ�K'Wٱ#&�L%�q�OLA�c�+>
?F�)_x'�y�_v���wm<u J���9#A��M��Oa��ĭdG��Dh]�%����e��X�`�Vxf|�u;����2f��2lw}'����B���M����(9�����q�������:(n����+�KU����l�
�r��s>�$��i<�M��$QI]�����M�y���8��h1:����R)�X^�b��L%�[��g�U�ev�t��_�8Y�4�B6׌	Oˑ�ңx�	J��2BQ1��J~�ءov	�ԽZͲg��lPM���9B�B�����`�C��~�=ɛ���줿�:K�s�c�ȴ������؅�W�X��)�(R�$1��\�js���UV���é│Qu��Q}����#�G�C�!�?;�Sj�02���F6s$$'g^��V�G&1��Mo����У{���!F����1,����5�F[�)�t�y�E����.ځ�A��CM�o�xЍ"�7��pY�߇�0�gq���A.�<6<,�9�|k4+"��OD�wj��7g���ң�F�t.dH9e]}����{�3��跣��h��Ɓ�>'Xb ������|������/%��4�iSsA-���z#��?�I5XMPOh|�C�[����6��� �)LU���ݼ/�}Qh��:,�������m���ǁ���X��@�#��yRJ%��l{�E6��N�a;"H�NdC���rN��6��ޙ� 5�
��ȥ��$+z�wcDȬ�Y'���y�������4�Hx��1!�:J9�\\�P �;F��ѝ@��2�i꡼?j�M�ꁞrM��Hϗ�T�|�U�^7k���������3.�+Ќ���=�i��h���L��	��T�����n�	�M��O��o��N>��̶��LD����H`�q��	��u�ԟ�MP�g�?�������ӓ/��~�O�{Cz60=�a��-?�s����	3��8�C�۹E��گ;���
��|�_�&�l��7�!|��i��VM��2�'��,����Nz{�
�,�~?B]����N�{t��-Dw@�A�K��3�mk�Ug����/��;
��n�"�  ���1���'s��oh��I���_�;��̙}��p(���Y=W���Wmfs``A�d��?ЖU���
�F�ii�%�:����ˢ���FEoުL���F�ײ�&�u"X��n���U'+���� ����K3  �֬T�a�d#l�e�WagI�zt]����͜���Д\�d�&��Lu�Qɍ��GU��[����]��ƀa�s��D���q�ۘs.�gF�J�?�qr) rO��1'F��ĥ�`A�h X5./��?p쑁|�e�[���e<a<�����m�M��M���l�{��,}7ٟ�A� ���o�/��s�$�S�f	��`���c����M&������]iei�X��\��^���1F�j�n#If����M��PLoT:����F1�����i�sH���=I�k\�6UIQ�vIl��[O~���,ȃßEh��Z&�.H�pc�����M���MC'ʈ�zG}p�nW\�O0#��00��@J����(��n��Bh�[1A��n��B�[D}��y�~�G�����,πws��"Sr�HV���v�!���� �ط�/�Ǧ2���_�(�Fe�8�v�P�윪�m9��9ժ6iN"{���*ѥ��Sg~�Ԧ�O�����_��b���(��S�]�f��yáҏv�+���o������s<�P��{*�<�6Z��Sޯ��5O� �{�A41N�nx_�X�D��:�`�br�?fL��M:?�!u}�q�)���g�O%θ/�D�88�[�U�E�h�(��'�~n~��lo5pm-rc���������b��� ��B�qٷ��6��tv,s\�
O�J�Q��oWZ7���bhL��Rt�٢�,��z\$UԄ �0T��OJăy5R��p9�1��K<D� �c]mr�4����͛}z�c��Q�����yЇ2��T/��~�CW�Ӏ��qs8�4ΕB�����Ó�/�"�����BrҠt��A��m�Oq��j�}��zK���A��W�!�� ���+ݥ�j�!l��U�ܴ���xi`$S-+8s���)$0�_2�����󩺢�"����U"e~|G���ti�θ�u��-�F1� ��F:$hk��!.Zq�>_���׹�������?E�����e���}��L ����~����i/<���  �@��j�3��?�썢�p-�~�n��>L�����r���M,hk��8M�s���4�[�}���/v\|�n�K�v%�!W0��/�J�=�6�#�
�z=0E��N⫞�m��l ��<~�e�=����[��uy��7&���) ��;u��~�3�YdMH�yb�,����mM���Z����$��=3c��	_�E�B��l�`����C�K�NՑl|��R'���2OJ��|��_����s����i,�#�:`���Q�VI~���/mE~�~z��U�d3�;e�m�Ȍp��� ǩ9*^l��ԃ�,�H�r\�Rw�J�uv�-RӰ^�&6��"bP(ҝ�*i6�D?�^f�z*��E�V+�N��F�b5���t��I49�8^ͳ&��?��ֶzJB�(p�>����Q]�e��.�S:��41��>�����=�x��pG.E��m	�o��(O쪈�C�@PW:W�+��2R64 �@O�����L�ԖL[�Y�iy
�����u{�z��GN�t>{\J����)Fs,��<*��@��D� L1_`{יB�EJ' �N㓷�9��e���o3�nq��!�D�Ւ�	��;��Mփ���.����}�1��=<�չ3s/)
��ԎH�;�R�X���߈`�\��b�����<��LR<�ʺ"��o�Bo�/��@�[���h�k�_�R���<�ά��D�Y{�M����RB8����	s�H����w���ad,��f���� �Q2!~�@���1�p�Kz�r�FeA�"�6qx��MN~�r}�n���s�yد/�U@֑�v��L,��4����Oo͖�p�X��3�j�sEn�R32i�Ӣ�Hje�X�k-�,o�Hܗ���Y���=qNDP�r�RW`<+X7>�l��e�����	�̎�v�A�BwU� ���ȅ��6�{s�$��y�E�l��a`J�o~�&�<�%%a�K�V����q�LW���5����?��W,��,��0�n���y�;T�_��֋.�C�D'�;B4*Q���:���=�;�M�5�jE*������V��v����:��x�ʷ���ϸ�$��ڶ��G<>#�W�R��6����~�N�Z�d���_l��7��Ί����?����^7�Y��{4��C�/�v`��="x��d��\�g&w�J<��i�Z�M�lAby�����χ$���	{�L����c!�H�?M�p�S�C�l
��Ea*��`S$3Q67m&0��\���_
^0C��B�d�뻘������ǅ�����v:ι�ߧ�� k�R>��#��n|��>X!��Ɛ��ɣA�?���V�����#�W��Vz��2�^��(�yEw�1S^�"�!L��䈂�X����x�Ž�_%�!��c��^m�^2�(�BxA��[�n	]����b��W�>S��	4Hm"��L{�T$�II��x��V��	�5�4���&�lMF�V���Ҝ�%#����j��)�P�V�Tc��Up=��
U�s�&(����+��biWyV՛�� ^k�F���h֢x�N��o�qD�܏��M�+N�����x5Q����V�ȋ_̫8z>25�&�V�-M���7΁��꧜b� |�Q����Tw�"0E��dm4jn��g��xQ����;۪V��!v��:��|��IR���ճ����/w��&R� :�M$���>F��
μaLXAÁ`��t%�T�gF� b�=��� O7$I�C�K�|�K9��5�q�X���D��B�b���dwv���.�m*�G��&�B�I����%LQ�ޞ'���v�1�e]����պpK��]#*@F�P�qV\&W��&�Zg_��q�p�D�7���g0[o>|��ق0�h�K��B���+�ҋ�Ǜ�}�)�#R�zޙ#tCI����ԡ��T^�^��g�����+�iХ�������@�m��������+�m��]� *��?8[����B�46\�5h4�8KXC��7��IN2�uN��8��\f%������N0ijTt?4�:�!�=XQʔ8�����soe�����Y7��@K�2��ʜq�L?AbF^�َ�y+NU�<P��<DG@E�~PT=Y�S���g��nB����˯6�a��e�r�ڊPv����%w�<���nۋ�5<ͥ^͇|�^�n�Wrh�[/�ݖX:��tc�3�$��d����_R�I�3����2%�G�K�[V<�i����8' ����~@�cV���Y�Nu6L�}2׬��ʌ����������{Q��qn��g��םJ��5�S���2��Ye���
��9���쉯�V�ʜ����	a�;�����?]#P(��7쮛�`9�����|Zܣ�㊾�^0}C/J����9��(�>(|n	�x��{�䔶* L�^��ئ��GYn@"���)o{����|��5���~�{��z ���n����j��`�r>����vo��`�#ٛ8�z'����kED��Q:.��yeچ��+�v%h ֽ�@�\4<���j����癑���~��w�����m���D�2���:�6�(��L�Y�Eu����WE�᜿��%N�	R�k��[�e>lg[�!y�(����'�A"򠐦<Ä��v���ݜyHէy��l\�/�ǖ�ke����F��8�EGg���nUQ�r�em����]�V%�o����0�j	ʹ��=rA�pR	�ۤ`��3�;"'�9���O,�jԄ���T���Q��1�O�4B8r��TW�ht�=Q��}�"(e�6���m���l�
��K���)fk�ш$31;�����nmIfsν�1	t@�l�zjyG��x��o���Ǯd��
^"��h�1l-,��t���~$xq���2����%��� �����܏i@�b�F� �����Ob�������xW#.ҟ�>�an[Ϯ<��{M�ߕNec�e�a�p�a Z����x|ܐ[d9fg�_{���2�\���D_��*9>��9�8��d?��>M�Hؾ2�@��)����8��+��6��^@���z��v���v8�z�'qǗ=K��<�{z�����ԜbL�u~���%�iO�T	C;,0�n�ڤ�^���$5�ʍ=����hxhh2�ɆW�^d�1�9��]EX8���΋z�-�ˡ[���I�M��=�NhJ���*zX%9@��s�����(:��!t�1ǏVbB��nܠ�g��2O��.�
�,l*�'��� >^�A�4�p9Cʆp](�>T��ky.4(ꒉ�P���s��/�4�n>�dX,�/�4���u������DF?=�퀄����!� dw/�j,_T��*�'�+U��қ��RZ��%���73�)`%mS�#����e�Ց�S'=�rR�!^��k]��:��|�ѕ�Ph̄m6����f�\yy�������`�W��uט�4a�k���닣 �L���T�e@�V��RKG�fK���t�	�4�0��i�5Ǳ��$tu3���0�4J[��oXަ�
�e�؎k���^}�`ƙ,q&|�D�B�\Y���@�,�u�S�,�j)��y�m\ś�]kJ �?�m(_��n׃�[���)�f��v���v6�g�쇀B���%_����0|>�L��z�w����横(c+.\�����Ӧ*�2Ո�J�hف�g	U<g�w�T�Ϳ<:�O&#:�d�,���.>H#���8k���_������L���g��7�tA�X#���~&�1%�o�[�z2����G`t,0y��������)<L"�9�ջ�)���h!K�G��pa�5�|2U�Y��cPk��������*�d@�ձhk�UY���cz��r��q0�@(�����kq]�v��O~��s��(��� ����X�q��i<wz]�h_]y�X�cpO3�k�5'��g.���F�C������y?8�����r����*�y���Y;G��\�������j"
.R4ޏ4���!�#��eu��	�*�55�e�X���P����2!AS��?N^<���eO�@d�M�%�.W�J��W�(��N���	xVM�%t���)%��o f����C��|�fF�Q�iB�k-q�M9��ڱD�$�8��9C�MH��S�#�_rv/�]Z�[�����vNX�X.�8�<�쨽3\hH���˥i!��A�GWT���ƽ'�[=ڋh�t� NLN��H��Z�sPDE��{tP�1 � 3@E٥�ߢW�����D��k:�mq��¾Gc^.�.UC��R�_Yͯ���	���qR�.S���g�>+�����|�p��E&���4P0Or�[#�?eḧ́�a�; �M,q����p��2�v�2�d(�7�$s'����c����f���V�����@�s�2�#dȆ�H��us7���6��=P�����!XV�"���Ωӿ.G��ٱ�]�3�3@�v�vǒc"��!}YQA �?Ma�{J$H��!�Q@lZfI�Ae��m��Μ��d�ѥ���vP���eP�s����9�Y�g)v˒6�a�-�R|���c�lM�y�P@�1������bl>��'D�^c�	x�B���U
�K�Ῑ�?����JN���3`�#kg�zL�����b��v�8v�"���/��n��n�*�T�#�����ѐT�i`��\�<����I�a7�ࡒ�\{#�.&r�����;ӑp�~���YU8�H�2p�棽����kJ6�s�A'��0�$��i�#�㧣��1�m��<��xni��m�)�1�;�9d�ɜ�s��r�U&����h��G)�(�(G�W!�,T�Tvk'��"�2�fq�	��+l������ӷ���"d�ٝU+��F�J2V�o)\ApђCr5�g��n�PErs��ÓA�����W�lw~��MsD��^�*���h�nU�L���K���zT����Z� �l��V�f�\��}�q-3�#j"/��-ɗ�G��e>�G�F
�]�,��zE�Eْ���A��~�"�aD��YB�4��"�#�\���bD5�%�^	2>ʕ���T�U8ٌ<-���5���4��C���"tc���������A�������2o�u׼!���#��zᔚUT���*�o1�?��i�����FC�xU�z�n_5��6v	�V�Z���� cG�bS�`��� ��/�bG-+ϩ��!��u.��1���6ԉ�(ZDU�ڑ.w�ޘ�7�t=�}̟���Sl`��{Y�P�Sx�ft���c�%�㹓%����Y�3�����}	�N���F��*LV�t����P\�ݝ�RE��� � �墙}�kT=���g�Mf�w��%
3i�jS�JENY�7k}��)��!I��U'AT#��7���Ǫ:Y��oo/����AVȮ!F����H`v�Z�/0|�����h<K�<��pm��k��Ma��"v�%������̥0!��KjrP�$x�!z��W�h���ts]QMm�:��ޫ���C�^�H'G�z3R	H�`@ H�"U�"�bhҤ���T�ß ϸ��}�/w�1�v�Xsf���Y���P�F[W���2�ǔ^�Z���\
�p�.�M�W�Pt#tc���oJs
H�h�~��_4/���d�$ጦd�{��U��Q�;Ls�kȭ�r�TD��+ݐ�xQ��*7�	U���Y�7{~7� ~�kW!����o��F�����	�X������_�\�wGI!=+�DbSV�z���	n�qv�Ȍ^�8C���{0�m$t����US�Ϭ�@���]�V��s.n�)=����(DM`�B����r���圏�?l�Wx?V��P1Ԉy�#3\|��J��W%yln���뱫9tJ_K��Qyc��ܣ�V��Z�[��z�HV����_П��"4�x2W:$�,��L�g�k�?��bec�΍̌�'��)'�]�5�6ޟ:�<@��\�A��'���r�
�<Nn~�Q��=���dM���X���8=ʨ���Hb�PzXU�d�/���m��a�%𫔘�c�VD\����L+�������1�����	\�����yx62J��Jw��O%�&u�1Tr;HCQj?`����D�@�:�S�h�:������Š�r�+w���1n���:'��i[�����aNJ�*�������ɞ�4>�����v�H��O��-�]F��df.a���U�bl:��x�Gߙd%�s��\&JΆ����Ц��)�X�@��'���\�1J��ХX9��mp(�W�0��Q� �i1�(���%kY�ύ��������b�Z�`��
<X���=�ʮ�h����71��ϰ1���}�{B�}��[b&]~`���Z�Me�����Ҽ�B_X����T����\_��u�0�n���|�s
��/����g��~����L�x�%�v�ZW�%a6����� �iW��U����Y����vX󥒚�A���'��m���k���7��/z�I�,�eݺ��'�#`��-��u(�Cv�4�d죉�+���,�z7�T����#�L>$��@
�9\�q�M���Mkߊ��jwY�|A��Qq�T��,f��s�H��Q�d_�Un.WϦ�3���ͫ������7TL����{ʾ���xE3<�+DY~9�%�DYp*��L���0��T���Adxs�9�e�G3��������
�m䲬^)�-ʆ��BZXU��]&T�K��!����;��5�F�q��SX"Yֱ�$����~�k���D���Hz�M��&+�nN�Z��)
��~V�m3����,Ӯ8)M�{�@�X�JZ��1�/�ʰ���8�������wՅzW��q����u��1&�J^�2xPqX��{��� ���D5��}��_Ĵ�6A����Z�
u)�[rJhA�5��N�n�s�.��ԉ�c�c� e��}��|�� [�t��P->ͼ1��Aw���I|�n�K����qJ����B�t}5z�&R9�y���/B�NIA� �8M�e��]}E}��u�1��R=�G���"�M�w��'�(�#�sOoT>��_���4d5�9ړT�ǚT������>=�����v�:�����Gđ&��`׸	۾9��Y�,`��]�2F�ݺ��S@Ž����y��) �')�{�=�A�9�� ��bL�0)�|�-��SzO�@���S ����Ŧ�����kǵ�,/pN@�L�GN��>_(�U��
ql�KP:�^:i��'@�D�hg��:$�yk�ME�p|f���CzzB7���M�2%`�Ԣ�#)���O\���Y6�j��,�P���	Bl�3�q]�=#PIj��d�h��ƹ>�����'�?�dlsv?�����ĸ���e8�j�b��<w��UDE�6�9!��x��Q&��eg>+ �N9��wc�ዳ7�f�D����]]��G��ô���`�W��}Ñ��Z�ޱ�^N�Yd<�Ĭ-a�{�(�
�^�/1AeŨ�lx�]���H���1+|�O�������'5$W������nk����a��K*l����.�Vŕ�Sr}+X�{�	�Ͷ���4<�Q}Z�x�8!K#��S0���܅f��c�H��zJ�
OF����������>��/�%Wt=�Ό��.��+&�ܲ4��Q2ҫf���`�j�ϻ3]���'P�;=b���D��ķ��U�Q�f�����t�<���.��[�F{��r����>�4�� ��u�>R뗃�/�:x��>�A|<��S�*'�a����Y2�v]6�$���cJ�\Ѹ`ѷl/���]��q��:���-�+}��տF���T;� ��]j�yc��~<3^�c\ÉrP�J���Y_�f�*b)��?�M�8	&ｓdZ�Ԏ�����/�T�$co2�ʌ<�m-�f>��\��]qJ���*f��&b<}J��㬷����ˎt����__T<۠�U��*�NT=� TʞC�ޓn��l!�*��y�GOYd�x��xݺ!q~蛫�R��=���Ia�̒����l#�ΔDj��fLXr�����,���n�'+���G�|���ؚ�z6I!�H ��K��V�fS�h�- �ӉCf�\�ޢ��vyO^����ٴJqyerq�N����͉�9�%�����_�2����%[��'f�y��A�Cm�.����[T�����Z&8�	K��	N�|y��6�W] O�3���1�H�|��?5I3�v=***�t?!�]��������&���ϛ�0\ک{[�b���X*(�ڦ*h岛��w�0k���S%�� vl-�#DB��_�41�텉��$���3���K_l^��6���%��h�ϫqֻ�^>fG��KV�_���"TuT,B�N�]�K7/`�.u}(T��m/l�qo��^ o�.��`��^g�) x��B^�?_�Wp�>��s(����[�Ǟ�Qc�p�C�E����V�}:�*��&�%���y]1t#�j�*,�:J=dS���b>0�:i�/����i2�!L� t�3���#�N�T�z_�Bz�y�ʎ�������mG�=���f��B��fk�kjǵ1��}���3���u���UZwq7���.���.#Q�С)��x�o�f&p� �@���F�HL�d9�څ�������)�u
 ~�jA`* ��ջ�zp?Hݢ�����n���(׻į>��Ҥ��E����z��Gk��ydy�k�1��3;V7{�����/+I�� ���7��h��>7/�r�
(�휥�L�bcc�<��aa���}$��s�����u���	Z��6��tVoF-y�1���xw$�g��V�����K��&���ד�dޞI{d�`��x8�G��3��'��-z�!�|����,��W�
�y�*�Q�����5������*���
]^6�����!~� =�D���u�$�u���CpP�)��v9�����j��Z}�����YJ1�H�Y��m��W(1� n��S@H��P�ޚNǷ4�EV�8\�l�~~Op$��]6��ܸ�lS�Zt��R�(��d�V���E}�����.*_�;z�I�)���ӱ���u��P�ym�P��_�����t��@�)�lI���o������k�R"h�, #�7yIu�`y��H������0�S���=g�Ȟ1�L?
V%����H��s���j�B��*����+g=��fo�������v��9[�K�ɾMG�����K��d�;���u�:������G�].������P @����4�Zt���4tf�i):���8`�C^��u�8���sN^����M�U��}-���͐���t��C��=HK�h��}n�3���pq�qU{��x���I��Q#�\����-|2N{��W�5A�)q���|�I��yC��I�Î"_�b��C�ly��ê���,i���ss����d��®��0.v���a��C�J�5���;�N*y� �ڕK*��Jv=�S �����o� ֟@�:�H`�{b�c��|����;>�D�^�^h��}�d���6&�y���g?pv>��j�8Z���Rw���­>��E��h��m�]������,�C}A�Uy0�1�р_ ��1x�г�lW[��F���A�]N-��+d���ޓ��w$�+n�*o��b�3;eBkU/\����"�������������/RU��X����;��ˮC���M�;ϥ?�F��*��Иn�:F~�	�K;{�*�Aq�b�W��j-�PL4iq�R�X*���C��ᮒP��<'O1�:[3�ϑ���B�ǅ}5W��AP���:��|����]��]� P�n*#7���p�F�`�)�(ؘ�	��1ơ��v����sP�"ȸ<T��ު��[0�+&|ӥ��Es�A�Ed�����}�qf��W��u#��|�y,iy}�ɪ��o�pR��%�E����i�'����9IY��P�_��ui2	���ߐ�۝(�w�O	�dR6���_�m=�t\��A�_kO�y-�R��<���֥>Dj7�1�R�d(�"0p�� ��S�:p�2�8c�|Q<�a#)�ެ�M�9xm��K2��Rnn�}u��
�n{�f�,�X,�)ML�p2�Itd�D��IW�$��;Bg����'s,Q�����'AJ��X�(�R�(��e����#Nm호�S��5���J�0"�n��5�9�F/���~�7�+��yG�gO#��[Q���6h��ݞ�>�~1X�	]?tD#��KK����Hk��������O￤e�4nl�,s0����ߥk�=��׀�0�������	gg��(z-Z����"&c���_f"��ݧ3�PK   �D�XYY5dl It /   images/1f408b97-f73f-448b-bb6a-3763ceb62f06.pngT�T�Q�7���� �HKJIwwH�HH#94JJ�Н"��!���]C�k��}����k��s�s����焨(Ic��#  `��H�!  �!  ^��^)���B�!�㄀�D����;yx��YR�����3����X�Y;��0c�w��z"@��@� +!��v�r�b��q~:p ���Y��FEUT9&�T[���ņ��*	���)�xP�|͚���*�y$���7S15o_!ll�����n�1�.�A`�iu�C4�(��������F��^��z�G����t
\��}G� I��u�)3���f��Fk���w�)E	��[�D�����~*�~#�ߘ���f]� (�?�֊A�#��GRs10%�!����*u+w���:�A
���	G�ϱ)|��|c�"�X�X�}F���=�a���@�?���3�������#)ٜ�U��#�L�P�NnǄ�/SZ�4I˸6�ʐ�1C8�W��$�}S��B��G&h���ȓKWi��ddy�,?O=g�P���ϝ��3k���:ۉ�_w��7'4���%��m^:9��X�Ś[Og����vR��y~9<�S��yw���;#��j=���G��e������1w�7U�C[�Z���J`p��4z�L���H~�X:h�,\��G�o�����7�׃#`�~������o���"������3�h�gn�!�ijD��pO���y}Ř�7�>����4�^:p���P:G����4T>�f�?�1�ʚ����?���9�,7�-�����=zU	=ť�.F��X��8Zq�ja(%����\�YJi��a3?��ȬaJ�I%�E.�TRk=�݄ט�%U��,G۱ʪ��i���y��Q����I���@��{Yb�b���[��DԘ�G���;~}(��oZ��ˆ}��v���uDPk��Q&���y��R/��+!I��lxB�X���G�n׶[���>��k���Чͧ�O�Æ���x_}�V>'����ӄ8C�����+��6њ�XSNy�bnWZ�|�����F+Ҳ'0}h�bU��Ἳ�~�w-�=��x߆\�*�ڷe��]q��5�5(�M|�.�|k�qڀ���֢ŅѧTo�
�K��`��wR�R_c��w۹��d�t6�.��)��K��2�������/SG�%F��m�ꌄm�r�7c^�7p�0�$0� :� Ю)�,3�Bkj����3�� n�LY�K���K���[��z����Ѹ)��~o:lE�{�3�?�[�u��W��(MV��H�utZYN�u��ǘ��o���|��W�%$���餷�V[|M��࡜:!s����	 ��[ ]$�2�NM�Z��JN�EA�-)︟.�v_��[/.ǭv�! ���SR�1�-������f^b	�oɖgPu+㖨w��Tye�Aª�7;"7^=����@�B44R�u�Qxa�8���#�H��O��> _��V9g�����fJdq؏��"��#����a�}1�G)Z���P���	̲��jm����g�? X�ӑjG�XZ��܁$��om:��&c��'���
'�B��k菼a�.�tJ���U�:cy46���������C1E�V:BX^�^���X�,�r6 >x|*g��c��oN��>�j��V�Ί������Z�K�v~��_���ؿ�/�eց쉔2��n�E��s���fk��<�o�6k���RZ��!�[�5�Zn)w�0�iy���K�.����1YJә���rmo�0���܎ޣ98Hx_�<����M*U��}����Tmoo�'t�_ڪ�[xE�p?��}�yA˻�U�g	������*D�	����%������l�u��X/7w��1��̛*/e:�/��7y�L��c����\G�<��C�۰
Y��T1���${:���B-��  ���*���|L����vY�Nc1n�Os�����6����U����q���O,��S.Mz���x�ǭ�rњB��/eZ�+���	YN�:e˺w"z:+��?1OF�訣9�_Dh��]@�{��A�0v_bP��=�x�:BO�Qx�C�?r,g��W��c,/�3G��&�P*B;6�+�p��?G?n�q�_}��m�-7��CG�xM�x^�����YPѯ��+QթG�ݐ��dE�ߚ#�i�o���obN[�z��˷QQ:��ΈC�wMM��R{6;k����������G#"���?�o�[��F֐@�����+`���%�v�}5���F������b�08�NE��43W;��4�_�89Yf�$v�M�5r�����7�J.�B�)�4�]9��b��!盂-�����^U蟫�8%��._��\Ƕ��a�����:f�V2@�)���X�X8��E����c��YrҪ2?/��r̴LWr=�B�IΊ�C�t.��{�Xڹp)�(2�y�����`�3��~���cG�6}G�����/wMF@6�A�,�
�ۈ;2ӽ�T��9��xQ�X�Ե)(�n�r��~�V.90�;]��+}x�e9�Q#-�
�:P7��|~�l�b�.0o� \6�R�4t�>�����A�Ygk�	�u��
�l͍	2'QH&V��bk�1��B=t7pw��x%���Ô���2�tS��C�o�j���P˲����nZ%j`|U��Q�	`�8���X�I�o�������[��T�"%#ٷƏ�eRpŕ�o�)tn!��b �Opk��*�Av=���R])V)�]�+��(]�afx�d��"cK-x��\U��������A��#�W��7�Pz���,Z߃$ �6k�CXX��;
$�y^}���s�V�����q����Zo��7���	�������V,���`c3�Saɾeb��HFJ?�L��:���U�Lz���W�I�"�6PJg(:}''x��5��w���z7K�9K�H�[�:�3�����k����tY����۝�s��9�k$r�!D�'�q��e�ne�u���6�3�_��͉���s�a3l<��M�������

�v�~@���z8�%����<�Ҁ3���۷4p��>Ē�a�i�_�-ͯ&V����D�}{^@�9o��:�p�|x��;������1�#�?!��/���,�`G����4""�e�^^�&)eJAZx���Γ�j���BOL�Bm>k��|3V���Ǿ�"��<��0�r%m��\�Pv�c,��5�d�LV�~����b�Un����k>��p���M����U�v�n�����N�b��7U%���s��貄��cH� (�߽l�9>>�M7-���%���v3@1%�(�M�kQl��x��R�Έh��j���;&�9ߏc�ʚ�o�DcI�y �Ď����� �U��ܜ;u(��s�S���쨼���Y���I��b,�ž�t���[��x�G��{����-+�	�Z�V��t2|��9�K���H>�_��Ǻ����&�&Q8^��]y���S���XzGR�Q,�>p�-H R�s�� Po���b�uՙ��f��c;j&�'|Y�I��|���v~z�D�#����oD���Nb8ER$���(���j��5>�I��DM�,G�I����'��
�9�D�Jw��y�;$�st�%<����������U�<��]`09����>��|�<�+E�Q��A1��=�<17��۽��?�Бz�о]�b��H���a��P��!W�T�% T�˝~s����ا@'ѵ��!4�5�o	�TkM�g��y-�AQ9��*p�I�NR�x�?8}����8�A&g$��Q����(=x�ϙ�9"/�m�W�~G8��h$��U���߻�>Cf��_&���Mm�¾�1!Hb���!V�X��g��H�]^0�䭖$����o�a'͌��L��z�|��FlĒ>�c2:��V���� ��8 �s�����9~Xu\�x���N2�C�h��e>���ʛKC��#��ʱ�>���+�)):��:0�y��g�Ar�a:�,	����k�����L��(��s���=�ؠ6f����6�Y�]D% ze�K��+�$=5؋U��YhZA����t�ZsL �Aml_A�8�-�����q��������i�6����4AѪ��A��E�:_kX��=��PGT�}�R�j�/o���1K�B� ��gT����dh��0���ռM�H�ȇg믕����B��39��4�:]8-+�={^G��go�QY��UU��R�]i��o�mw��!R8�E��^�=�]�W�r^�@�zF�:�j^6&���`��/�	�*?|=�Xrų'h�ՒӜc�᧽��d#�j�l'�k�����1�nb����{x��ŕ�#�\����>�����ٯEt,RJЩaM�G6�C$�fm�.څ�󁃀Օ8P��#��,����L���.�m}m��)��������	�,A��f<]�{Q�/�KӁ�uq�Ԗi6c�ĉBi�Cm�o�4���<�TMKu6]W�&zaW�a�N\0��xO�����	_4�P�>�zc��19l�TS ��=>+X1E��ev��&1����y'h�է���V�����~�<g{>hy{X��͖)Ȉ{�~^���BYq�ݴ��Lx�B����hI�w��;���ߦ�cV���w��s�pk�К��2����#턮*�vS��p' ٱζX=�ƽ(Ͱʷ��%�(�.b_�)��n�`/��W���SV�|.��3�L�=K7�Z�}�x�V������j�� ���\l�=�߄�2 .� ;������g�Ä�D�r���{`��	sy��R'~��U�{���S�Z�l�M<�F�BTCE�?���qfk�!�7���hAqB	|��bN�Yq�E�wZ�7�A~,SB�VE�&�z뛍9mټN꩞�7v�¡\u�� >��4��y'�� ��G��fG	�e=�����׍i)����S�.+.����j��%�R44=�Z���,נ��ג�j��Z�Z��G�	1ų�]]��gn&�dK��M���=\��Y/�T�4�e.(xz����
���d�bhƩގ�KT�1׬V�:�Z逽��U��L匿�a6~8����h�߅-��@%�x7��� �*�;&(A��˝�+��ѳ��V�!$�����`���Q&f^�l�a��q�F��T<Y��L A�e�?����:D�Mđ"utC�
�$(�����vv�p�Q}�0���ӽ�R��r��9�B�qRQfF�W�?�}]�}�AY����G�i� ��;E<8�nz��'� ����P\���'����c'tY��h��lv����)�����m|'�L��%���銂��hJ���s'�C���u�� ��J���;�q�G<{W����Y���B%w�C+������;�;w�6{��iz̗Q��4�gi~64���q\T�>��G:JF���p ���^t�c��_�ԩ�
\�<i���}��K�Y��ê��@���*VÙ� �����~�7��?��Oz��s�й1�~|���nt��E�r ����UF@����
��x�"�(�{�ݗ	�*��z(2�����%8�C����pj`��6ib�U���2����aɐ�cV:T�3�<��яO�e"m���K[� ������̶(B�1pI�s����2g<	=!�G�{�y�^/���T�v<��Fx���دX�|��_��hxz�����'�=�,s���P?{h��T�&{�t!���t���⏮O�j��5���)����P�*[�}~0ELa��b �n4��I ����v�h	�gY�9�����l)m^z�DS����v?��F�cE7t�=�V���y���S]tI5q��2\ڗ<$��������l��>�,���W���m\���k�$���l�ph�]�3̙)*�y�ܜ{(�&�E	]x(@B�n-��tk:þ���r����0D�	E��B�.�V� ��e���J��%X�aNx���6�y�������A񅇛�����6����&u�^��C�ӯ��X�X��o/�c�BO� �ȂkA�GOJ];r�o�-�2�=�eƟ�  +�7=TYqxM��G7&g���~TUAQ��Wz�����0�g]���\�,�|��X���O�S��1����T9��"��[�V2�х�|�/>�Ԙ��x;%������|!��{��EqN�g�հ�P����;�2̗)ǋ�������i����lHt�	<uc��>n��L���D��| �k��ßN@J'�;���,�FR�O����:m���(d�/>���n�_	��2eL����O���<tr��,	)�ߎ�C\��������\	x��C4@:i�/4.y�lG�����	z2��{īg��E&r���q"w�RS��
�'$�.�L�`>�^iU�����F�����1�c��G�3���~ĸj.�@``駟s��7'�*�m7)�U�\o��l9�i��$����9ߣ��5���"?��%_�R:�[g��u�M�Nb~�Q�7Fq�?g$u��r-'��,!*ܖb����Sc./��^%)�o,u�ba<& ��(P��m%2���ב 5n��n���\��2�&`�ZL,��D۳�Ȉ�A�1f}��u�[^���,vxn��12ܓ�ԤxF՗���z���_�=zm����h��><��b�f�I/���Z���%l߫O�����;�6mmc�Z.7��x�g�ru;����h�,��ɍ#����T�ݏ�pʂ�sZ`���ج�$�ј�e���c�)^�� �LV�L��XV�p�&�=ϯM�b���?��ay�m��Q�!����:���]�d����n��`�w-wŢ����׾%���i|ŝ �U��>��4ٙ&� �T)���[ݖ�z�n�0ǉ�n��cm��Y�-�WS�3����ZJ�q���+�'�4���E;q�b�c�pH�i����p�����a{��(�킞��ť8>Y$3]�ˡ��:��Bm3IX�l�M����|��T��nM�0��6�>ű?�L� 1`��T�:�w�k�V�7�!u��c�>{*�#)�0�Z����;�Ù�;��Qmo�[{1eu!7B���lJ8v�\��e�[�X�w�l[ �Y���S�AB��`R��x ��xF�Bz��-_1��Kxxg�f�z�7¤'�R:�(ꟶ kx������U˯d�x@����<��
?�XS�H�3���LL�)�]@�8��.1��1Oi���m���_5`q���z�l>�~�6�iZ�Q}
<BK��?k���O��v�����˛�����z,�@ ]���Z.t�l����\�P��8@�������kU�=?�����*�����2��vM=�]},�X��N\�X�������-ތ�n<`).*$'1���E`I�>J����Q@����,��ɷ�UCi������4����9vF����y�Kuk)���G���}�<^�x�]o�^�]��Gu���r� P������t֦6�2�����$������|o�����#���L��8���1�uu�M���-��%����� 	l�u�,���a��o��I�r?���'���W�Q��]�j#���U�9�nPI�aez���	O%�*+����z�>��	��?]L�:��/���=�>�}����?Z$J ]ނ�\��3�4�bn0�כ}�b ]��b�;��[��FV��s�Xq�0�N���j���u� }��u�kru=^���3�F�V���	�p��ׇҀ�F���Y����"I��ܔ�!�#�\Z_O,m�dkK���P��ԧ�w3�)�{���[Yet�5�H~��+�,�r�Gh�󟬂i���<F�/t�l5F�|~Ȍ���U�Q>4��#��̃sn�*{���bT�W&-Hz,�z�����b��<Kr�s�J�����~MFx�����Li�yx�A�s��V$�N��v�-r�R��GF(�?V诣��۴�(s5�����a�	$54�|��O��-����?gJ���G��"^�[b����2��d����0� R=pn8�0�ݍ��ʾPc�ӧ�FO��9�r!�w��|����V�-����S#튯�����Ś�ߞ��l>���B8W*"GK���������	*�g�28;�%��vb� �E��׵Ī#j~C;譀{�^?��<0P@I�Lj��b��h@�W���I���\��x�w�Z��SG����/|n�_�|����j���p��_Nu�@�N*� �>,�뿽R��%�7����5nN,D�؊L�Od��Bk\�h��"	S�H�v�E{A��H�4�ʃO;Ď�"^N�VT��`���V�J෺���i�V��%}^�~MkL������Rq3w�����G�}Y�34Tx��p;s�u]�ͯ_�|F�9_�.�涁�h�� @�xYB
_��v$��W�/�X#�4{�}Q��ӀlE�S�-rIC>6��(�^�6�g�:oc~8S�xX�u������k����pӽ�lj::��%^�`��4o��w���~���*���z��L?��ӫ9s��^!8�F���5�:Ig����G�?��k�nx
�ǟ���i����D��.�X��v�K<��v���h����}g8� /Ҍ��#kQ\�]�j@[ֱ���ɯ)�|��T��}2�'�/n�.T��Q*QGvƑ�¨azr���z��Ţ,"�I��4y�絛�(��K�L	��� j�$9y48�:>�����V���P'�uqsZ>��{��?���($���u-WNR�o���b�V��/�.h�y��^5�0S�W9�!d��Qc�;6<���/��D���ɬR��B��u�(S��wy,o��?E�0Y+!$�r$�W$'�ww*��є��������$�'B�b*���R��
9�;�BO�s۳8)���t�%׸�ҁ���[+�	n�a����Otl�5�l������ ��< �D=Z���5,>��p�
]�5j�)ѫ�����V7$2�|0�c8!G��[>������ �:>��P�Ѵ2�EYd~@Y�K�J�xCI��H�]�QSyp �g��BF�f�6��t��h�$���0�~��VP�l�V�;��@����rֺ�s L��â��g��u�i���#���[Wq�]9H�����z~�k���ٽ��E��OVʠ�N
*��>}z���:�;9Y~O���̏e񲔑R4qy+҇�_����V���/�n
UR%�x�� JN-��ʫ@Mu
�W^ME���aDC˘�����sIm�|���즨����ܳ7G� �����GG�����x�@m�����q����a�� X4�R�91�ʲ<㔏�h�]U�u�o����7���;}7��3J�*���dd����'Z�(���؀P�2�������mR��D���=^p�f���(�vA��r�p�U=��\��v�<D&�x���$��9�6�8{�	>Et���Mx�d�'x�I�P�[��`�6R�n)^�f�7v2��PӰ�%�f������/��em0؋$��G���R���Q�]����v��D�CW��oK��D�a��mw�0���-���ɭȱ��w�YNq�Dg���GP��_F�+s�f�sb�*HlxJ1���4�4>�������`�[�!G�Z���������0��
��~G@��m�j���6r'��砥��O�<�ܡ��b\���j�>�ەk�ݖ5�_�U�u.�6��O�)P�bk��c�v�=<'���:�*�Eʨɣ�0?5l�F=OkŪ���eg��҃@ ��8��{��J�O�͓�ј+(qȱڞ}��o_�|&��p���vpp� 勓� �](�]j������I�*潵�ȑb>����'���鍥%����m�pSvcB�)? H���e���qYHp��D��_O</m�A0���+�2���(5��_���Q>��9��>/`��h2Zϖ�/Զ��D�ZK�����*�g�bM��$�LZ�'���R�����E�3 ���ߵ�U��Mz���nA�L��R��Ϛ"�*��	yk���T�^SSi����	ɛt7�����ǫ/����K���9lx��~Ne���q����(�؛O���p���F'S����ϒ_):�����b��� �+�~8�����wx��,A�_��d�f��x1���ϣbVa�h��'�<Z',cm�nt�Ai6�,����F/M��f�[e����^$�����w�u�FL�,�=j�h�/��?�rv&dF�ϮUJ���U}b" �jV�j���`�vk�w����@Q��7�-y?�åg�ӥ����oJΫ��z~��g;���z�I������B�	�M&��u8����M��8��b��2����#j����+oA��ի�x��dm�{E��r{"�j�g�/ޮ(ʣ���;Ȗ�ޮx��.7�mj�����ğ��t����$�_W�d�+#��j|��u�W�OWF�P�Ϸ-�]k�����dgeu�f��( �)�_iy�,�+���7Y�D��ş���1	�N������6[��} �3�V�9v6S��.������G�r&���<�cj���9�4�i�5'���rJ��2���$�eW ��˚m=�� ��=^����z�0�\zzj1K�O�����N�x�ѡy����c2e`�9�A^q|mK��D�����Q5�qw=�^Xm�ޢ�O`Dm�%��%��.�� {��?B�^d�l��Q���s�%Lm9I��7�R������_�]�G��z6�f�c�p�ge��|�A�F��s�LkM��m�BU���+-C�i�좳5V���mb���K�&l`V��^"���m�+ WNÏ�?�Q��ܐ�f�D�;�hgi�|9ƲI�&�I�}����(��/�#�!ӥ�(� ��#2�1�J��]Y$o��S����n;�h�QTx����V�I�2\��u���	�q�ֆ�
y�3?E�v�S["8���N��W [��G�������#��m+��ŷzBC�[߼�ͦp��T�1���ܔI7`�P���u/������p�[g�hh7��?y�p\0��ɺʽ=_�5��Z��jp��S�}�E�no1��*B��-?��=o����yԅ���b
6��@h�h��	��Yor�Xn��^=�����ĀV�e�O���}������H`�@.ưa����si��yݚ����[#o.L#�yC��x-����}:�(� A�ȼ�M���'VmWk�/�Z7]~��3����ZXP�eڢ+���9��9������'���(d��>e��D3�_?
¤�_����{�y��sh���)^���SD��Q�a���$'FJf<��ﴝ\�4��!�%�"�x�5ޓ��aBg�˹�q������p����x�
�_���q������?��\�^Y�4�~�}�����$2��z�O�r.�'qqld(��#����g���xp'�r7�P���x��>vw���8 ��`����D�m���=�OR8�k ?�V��f�ί�6Q[~�m�!�ط�'�_s���X|||X�$�3��[��%&j�I��D�E#��KK��#I��(�}N�d���Ǆ�MQBM��0�'�����M�M���Ư:_�5GF��j#L[MM?2�U^u|b���!�d�ݒe'?���1zs�Ǫ/I�?戤�?��*U�6��d��Qz �*���/��q�����s���[��[��vQ��r���:>�+W�w�r2�Tx�k��{ϓ��!��Z;��`Я��(�G�!��Յ�[��}h��CR�׆���q�k+ ^����AO"��"��_�֠v�U ,�c=O��3�L �*��f��WrC->�WQ�*�_*>���E	�������^*i��@i���}� ���é[?Zٲ�^�t���h���6b
v�в'2��Þ軻~6Ds,77�*϶�B����!Y�k�� �N&sv�΢e00���e���Z�͐��WgY��h���T���FPN��B&�l�j�{n>IB�`by�q0�>�����b�+t�_iǋ��%VN�OP��I�L!���F"x�ji`��UF��T0��>_�����$C�m܍�
�iy+h,�}��'�p�TM9X�x��(Ԯ~�Ǿ�K]�Q�1$�ܶ���K	��q"�P������p�'���]�#������o=l[�Wo��Ҋ�J���1�A����O����s�<Z��C�d��e�*sfz�r����0IxMп\ٽ���:���o�	BjD�����.���1k��:��4y���MDz��xZ����y��'�Z{ב�'�7�4���%�,�3%L������>��X�f�=��߂�^طNWn���;���J�m�cћ�b��s�R˾����$58��>��a�i�7��/�Dk����#l8����ى�l�>g��d,nãi:��'�`O8o���}�щ���(�%���:��z�X9]��VG��q���ӾZy�����L_�6������L�1-����㾰�[��ܨ�����䎡����R���-n�<me�j7l�)do��Κ(*KOZ��\k��f�d1@Xe��%�/y��K�\����7/�U��N�ސ�{x+��n�M޵.k
��gN@��H�Z΋ow��<Z�	���;���P��nI{���`�Au����|h�]_��~���)'�e�u� i�y�ф���n���U3���M�,�~�-�,06���BLU?����Z�F����TO�;8�=�L���G�RL�WĘӶ!�Y���gԒ5��^m�"�<����d'�?��j`Z���:!���Y%%W���`2��v!Q샲�xF�m������)[_�F�?�&�31H���x'\�1^y$���Q+�0���=jv�Z��v��M�G��]R���Be*k���J�k'��*��}Խ�����W,��c�m>;BO$���E[=c/�gET�ʫ|��K����-����^�ū{�Bx��u���	��F����� ��'q2�Ul&�y��&�� y�PAMG,}n�RC=�L�����`�UE����=#R˙�H�®i�ֆ=����΄���n�#��)�(v����y��ذ^b��+p��i���)>0��ۉ�����#�/���a�A��zz����M�,[��Yǃ��ʋ��c�>3%v��q�RZu�����Z�nd��1�����	��}c�4f���B6ּ�ULvv�M��o���Ͼ'�^l�/�Зgd�3STf������~qI�ٙ/�ޞ�j:4O=�xy1&�`�s�da���gO�/�ކ���܉��5tlv��\3-w�Z�@�ëK�*k]���Ob���jѓ�^�<V*L;�uE��pؗ�Ҟ^\�@�ϰ��@�8�Q�l�(��x���ΊߍCi 3�_�P��4�}V��@19{�_�*��Jc�!1	�
������GV7抉_l�g*��PM{3��!$zF��]���Z��!0>���ɬ�j���1��L�խY߱��~����,ExZ� ��KaZ۫m�rZ@�����NIxr�9:�Y'2�}q$������C�e���qM�}=;Qc��`�0�>1�{���\\.5]�!!�����4����R�E�U�#,Xp�,.% ����֔q���7��|�ZZ�ҕU�ջ��IJ�]^;�Pc�K�Ԣ�hŋ�`��M�d��O�9\$x�gg��ʌ�[J�YQ���ߌ�����V��f�K�u(��-��W#����l4I�:�������L��T���z� ��oOYH���i3j9}f��"��R���	��B�ԅ0N��j�(d%�X �X��d�N���v��k�#�~�^v�S䗔�
[^O�4��匘/0��6�z�itEuG��=��qlF�������@]IU���u�t@�8~s y��i�\��Bڡ��bZj ?xX�e�n6���	Q���t����ccR���.��y��i7/6�'��+���W8��wU��%��h�'��PZ�)z��F�)�������O�����fs�C����T�c���4�1�Kh�d�u����Yq�e��[6�w8�<E&M'�k8����-���4�Te��"�a��qYpw�Q�#��Z:�]4�]�=�Ns���w)�бH� o��V߻��[���m\�ѣrQP����(���Zn:Ȧ�N��t�E�.4[�^�Xq-,�91��2���+��Cm���*7B/[��>��!q���̫?aX�ژ�y����?��9T_��e<��x�!����������_�d��V��"5�^�m�B<5� ڣ�=d����_I|LG�[��Ҭ� h����jE@]U5o4e�,"�WsŭHv������Gm �����.��"QFTe�}|��_�"��H@�9�-l�3�`L�颂��������v����P�lB)Dn���G*�)MοUq��XKF�	z��q�oǩ��st�8ᯩ_��5�x��������w3&N��%���;�ܢT ~��k2�4��&;�bTTЬB�XF	��N�Hu���͑e�T�?~�,�ʸS��&�-4��~ru�E��K������s����y7ə���Im=��{�<���i��RF�F#I��ދ~�p��Ӫ��DG�c7��krc�8��/*���۾�p�s�������[+��4dh{��7�t�+-Ƕ�^�M���`I?T�4�ZG@�u�����ˤ|�������]D���)i����K�rG�i��Ú����u.�]f���1�̔nk�3Mja�E��G�'�S[n��<�S��}{#�v&*��K��������}53�,5]��Z�K>�Ip5�Y�D��x�K���y��'RZr���e��?��[$��[V�A�
w��!j��2�m|�L�,��  ��F�'�h2���v���^���G�~˒��H�*`��,�oٌ�3�c���i��Cr[9eK]��@4��V}mg��V�+�O}}�͠��:{6z\��x�d�89���	��jN
׀�&�g��O��X
�%�2OC���{��A���}p�����y��[5[�BQ`$,F�Y�4��r
�@��Hh�:(6���<^<�^]I���ur�hH����,�t�*�{4[>�h�%x�(is����pE����!Q��#���QAN��$��z��v﯋go�3�Wb�0��W���~!Y��>K�T�%���Ng!�{��o���3�e���{O���ۿ�LD�� �[/F���Ϲ�iX`����f��3' l"vS�_�V��N4��J���i3)�	~'H�J��34X�i
������F�G��2[=���t�\/nN�lGI�h)+��S�d������fr���~�.�-'裸��MH�55�Рl���6�n��э��a(���?�Ft�׳��;D)�0�B��_����$U�aZF�G��ir9Y@���t�Ɋ
��G�<�������4��@d�0�L�y}r�p�%���f��}<�_2&ԝ����$��S�r��tH����r���Ώ���Ti`!)	�p�ʭEp���-�u�D����C�E�jWbZ��*1�*�i�s?���cŕ�_D�M��Ɔ	-�x���7W]?�f�}c̏1A@g��2隶��������c�&~ƚ�ȡ�U��JG���4/�떪VX���,Ji{�"�׽ev=�u�F>�O�x�D
GӅ=.᩟c��9�^T@OTj��ƨ����y�{�ݗo�n��|�A!����ȶU�L�%7*D�mX:
��1�Wp�/����N����&���G�����VV���0�@>Ϧ�ő,!���
�0����6��G&�#�_E5�>9@����͟�|Ed�Ý�!{2�,�'��p����x�ka�^���F�#���Tİ{�ݵ?�8��ˡ�/3�F܂$��c�I����?��/���!w����s�z�(�Q<uc趯lbBR���QS?��8Y��Y�]�U�E�`ۜ)�:Y� @5�d^����U7�� ˎVb̔�P�+S���Y��;��r@�����&���Dk:��xz��1�g@OM��[��>��6���|��;`|ԭo�R$�)��1���0ϋ7#'AFʟc�B�ӆ������m�������`r3��Vdd���|5�
�A�N�UB�s�)�O�8�e�n@�/7i��-0X�	�in=�&M�&� k�u>0���~�sN}�P���6y5�	`���F��t�;1��8�7�W) ����\��AU`o��I̷LQan]�D׫�J��^�������ܫ���s���q`���)���oҦ�1�\�	���I���|*%l�z��s	&�ea`��MK*}�<;N�<�O�ȫ rѧ�\��� 7JG�����>�Z�f��1'��C���_��yaw�U��H�r�{ �ҤH2��!V6��������Vg}��<�?����ւ׹FnNh�sϻ���&CοsŧZkR�W�z3�����m���+*,�aқE�yFp2��|��:�\}A� ���"cq��J��b��2#a�����'?��^�zir�Pe@4��&�
M�gD�qYv�{�y�F���k�f~ƄĦ9W�������|�7�de�@u�j�*Ғ����+��xt{�d����0�ͻSR�OXDn��oZ�?Kc9�S4�m��$M֙�]�mZ\��K�⅊�4�唒?G�P����!��%pR�L{�\�YVr�h�L?؆�{Pݻ6e���0�.sZ��n�(�,�7�krw��U�H0�w�JWZ��I���7�t�֭օ�Iĩe`f���jp\�%����O�_�˥�(�C�t{Q1v�{��4�pW�N+�0�8�\z��w{�Zf�?��(���z����] 	����;�C�����������_�U�";�{o������/�Lu�mfNA��" R���H��d}N�|�
�j�q���?N�>����0�FU�9�OLx���ziJ	4���
H�IK��u�Ll�� �dܝHwa��X!��,�)w�W־\t�m����z����"7�6��M^��u腟���������t튷T�
�iB�oV��z��̽�G���d�\�
�C���b]������9��Au�b�`���x.�c ���C0o�O==.�*D'd߬��{��ۖ��u�$��]S}^��
V��+ܵ<m��c6=�&�|��I>��bg[g����MFH$%�n�:�a��Qm�� e�>�~�ۚ�i�v��JH�1V2�<:�{~_nF$���Ӄ
#���职:������'j�17�?��#�l�?��I1}���gӬq4�P�
H��k;�L�1�@�E> Y٧%-l]=ԯ�'�{?��µ�_��$d"�j���D��>>q$UR���`���6O�ĺ�s��q�a����&^*\V֬�L^Z[d=��!�.�%���1$��F4���(����Gxrf�H���2������}���60z"7N��4�vn Vn�˩�c��)D�ʟ׍8��4!	< 9BI��&j&w*��V��L�����X�3�6fJ��.�Nޅ�[�X�O�B��U8��jk鉬��/34��)�9P���r��~�+��ɻ�/�m���P�X�-5^���Oh�n9%�"��9��X:ԑ��;1$B.ja����K�#��\x�srFO���(�N��(�6?��6�d���P~���;W3����o6A�Q���kz����)�@B2��-V���SA�m ��_㜻�.z���v�oZh�MiO�_]�N̤�:�"�aJ�����(��^L�R���b�}�
������[�,���E�Eߏ��,V����O���+�#B�%��z�!�E�ݵ�E���ܐ�c�x�^�Sub��}�>�Rq�M�����y�P���W�?}�F�.���b��.{b^�F�����>/��yG��867�?'�ߛ�ep�*�1u�H���z�w�u���$����H;9q{_�4�$l�w�����;�Zwm�(�9�T��M��T-�Ta�[�|CMM�A+�o[�q~P��^^1�,E���t\��<V���W�3:(�,x�ͷ���-�ŭ��A��ܐU��iG�
��nn&���C ��!��t�uz�9���_�Y�~��H�W+�e&��R�}�l�����%�iU[�� M<J�?��=�w9��	O>�E�ƦĩA�T����0"�u�pT5CII	%t����E��ә[X�M|�];(iIK��߮���tLz��(�
#7\�}��3��5[/�V��0"��z�z��q�EIS�FOTCeTH®���-*���-I�wx�(�_굧�����~M��� 7L����|��e{�.�@�ō,���;j trrr �����+��e��9�+%t������ܛH�+�v|^�n�XX�_�܌�=/�n+FF�괏��0���^#X��O����gnR�M)Y����eH۷����A���7#�/B���*jjY99]HY4��y.N�ڥ��x�3[mE�|�#V��с&�I"����:�D�lTM��>ĻB����/�C ��/ۑX[gf�>	���V/FD{����d��I#�4_�6�N�X���t���d{����vy���d��i�!�F�[\�." EAK�G�����+h���6-O�-�S%�E5y*�d�1��**�D��Ax: ��ӉOϏ���6���� ��>Z��]% P�ѹ�7qrA@�(��x��*5�:�ʘ¨d#����S��\����Ŋ 	�_Ͼ�g�X�=A�%�#s�+�Oҡ�v���{�@��'��X�\���|D�<l�/����(nnn��_���� ~]�mi��Ss�����燛�a�Bu?__P�Ű�-����j���ww;�Wq'�
_�%� k���K�@��~��B�)�K��le���?��ު�}Lk������`���U:V$!��C��;� X=�'��o�闷�l��6�~a�%R�9�$7�?G���_�"��0`����e����S�%Qj>�P�]�Ö<DGG�Ϭ5��d�d|�?�;8H|-�櫦�5�-`�9 �t��+o�(�ϟ؆FF��0���:c�d/������W�m�����/�.GY��r��rL���X�¢J˺�f�[���WZִ)���;�~cu_�u �RT؈�:�wF������]���֖Gss�W4�]���� q:�>�jv>�Ld�t>SW�-�q>^--e���ͪ���ڠ��r����?���#Ý��H�a#6�u�>]/��RE��7VUMaIRo�w����s /Odfb�h�ʜtO'F���LKKC}\�ki�
�+s:��[`�(�1�"�,�5I�:����F^���O��/���<2��c�s����C=�����/lZ׮D244�v�=���ߘi�A�0\�����l���% ]tB��/�3|v�0ۃI����V���໋*ff�r������H����5��)r�jq�q��toİ.�T�j���#4b>���MD;�#�0��C��y7�����iİ�]��21�y���rP�D�j�8v�c`����mV�����/�))ě����D6R22p����qq�J�~�1� �+����QPP�V6D�0t&q���<c��ccz�|<gynV|DH,{�sqs�9��p�c �x���/�,�r��:C���4��7 PTOЌ / ���剫���X/" ��3����+������Ex|��I��V����
COO���̬s}�$(^�뿵�A�n[ld933�v5 �b�r��g!����HaF�I��Áœ�3���s�)�ߒ��ŝ_rz���S�@����3.HQK+,1��E�͍��p͗�VW\̲�*j{�z�q���7�z�%5�H��'�H�Oo��v�ڢ"�gA��ܻs=T�'�XdY�w� ��>�Y��I_��ߓ�SY�.j�a.e�\-}֌�L--/g��G#ikξ�s-d��-���'��w�5�s|��L�P>>H�O!RL�pp�H�cm�^��KK��h�������Jˤ��J+��m.PA�~��]��,u�AIs�'�^ꘇ1�m�N`LM��5}b�+#;�i������s��������7�q���.�q��9��v���f���=]4a0�;0rsa��ӌq�C	�<=���[P8a�~;�ySgώ�u��u]I����>pS����MM����8�2<�<���V/�*'W���v����w�M~x]��zީ�~H���Ě.����V�0�z!\c����P�@́�����6=$CYiU�\�B�i)[)���hlbbcj��k. �t��Ы��B�B�2�d^�`�������;{��m���a��h <$���Na�T+.N����'�*���5��-��:�l�򥊋<h%&Ko~�S٘��eVy8�� z����.OGP�4vDd!�6mt=N��v#��,]6���Sr0Ђ�V|��c[�ܛ���?�g����۟�O2~-&T�n��O���+���������u�-:��Q*�ѳs�Ξd2���+.n��>ZJ��L���Qm�{Z�P@��Q��#d�+��Wܫ#>"�'+o2l����v����˶�qY3�b���W�P:r�?>>��<{�
?(?�����d&����M�b��u'Յ͠����܂�����*L�?,�	к��`(C�[� �ӺXa&���j|���Y���\��&�{��VDY=����wFks��7���av��@��ۃv$��V�%d3��g��G6��?}��W\q�`���K��%�	t}�">$s�~(��$P��Y=���4wgW���,��n@��B���X�h��MY��8=݇�����1���l��.;%6G �!��\KT�@W-CC^�_h���؛O�
L�e�M�&Îzp�0P#�ȵ)����1��ԧ�Kt���ϱ�V/�4�]2Bw��L�:�Q****
���p���$�Ϛ�jѽ�?��)qÚ��\$�h����0���зg��С��Sf�a�bd@p��8�Ⱥ���
�~?�B|$)�ʗK&�l�ڃ�h�ϙx��|���)]ө��� �����Ɩ�ԥB:�z�4��w��+|&����|0�	ʯ�ع����yY������L�(V�).@}IG'�Gt�/�+�M��u���͒�0)��>�Y�u����P���c,	��� �NH�JH�����S�b�[��4!���4��3��cT�X����W�'�X�io�meMͧY��q>[� �uQ��9m݀��ȴ�0H��W�g���E�	%P`оMK�Դ[��I���e�R̻�I����AcN{�5J	�pAg*
?�u���|KUK��KW�0):l��j��
4R�G��\LJ��?������Yj�Oq:2��%h��C��`�ކ��Sq�`��-�&�����{���5Z��ߒ[h?�Yp�2q�>G��\��4Y��߰P�����F�	��&�w��a�*��mv���S��/�.0Q؃�k�`��#���W/�2���vD\���3�B&SB��$mmK�v*��2��1����V��tiD.���r�́��(��������MO[ �~��"�]q��[�X�����X˕f/	�7����b�O\�z����4ߣG�]3�3�"�1�[����@((Ϯ�x
1��}�������|�8XX
�n��b�%MM�����M��Eh�����M�i^�Wg=�'"@Eax��s���~((��"������zvf��Yw�X��!�fѵ^�݁�I8�f��pnq�ħ�����#���z�!!!a "#�V�vﬦ���ƛ~j���0O���@��)���d��C��[��yX@����fJ�CӺ#�����t�ə}<�Hta���̘2or�������T�8:���G�#��R��)�tR�G~�!A����4k�q4{HS�c9��F �`�M���ul���a000t�N��K�Nw�DԺ<��,0> ��X<��p��[P����f�F!Z����lyk�.5-���́���/���;*++�YYњ��n�N��N;j��3�#Ո�?�b��.�&���K�����
�3l~z�]Z΅7���F�D��z6|�F1K3�Q���Һ�|%X��mE~*�(PJ��T~�c�$��}���9>��ʡ&���m��r#�O�%N��@w��h��gEWઁv�	�ײ�^��$yv�P�~G�Y�H@Ǜ���EP]�sj���U���p��;;

��C�������2���1S)==
@�ޔY
�XA>$s4�[J�a�76��e[��p��v�o�ǭ�ܘaҫo�F�e�\(;�"��6������]�X�.9U'�����..F����!Sc��u��\��h��T�"DQVFݘ3ឭ=c���8�L+.�I߱!�tTcz{7��]l:��y8-C�12vy��Q�F{�p.�:A�����Vۅ$[>A"�������ɜ{P���(�@`Z��^�RH��q�,d��GGv`�6:))4 m�Ñ��1�����u�u`f�6Շ�x�F�����I�ǔ�V:G٠1R����qր���<����9&���R&.M�l����َr&w��;�C����8�"���o<
&&d��N"I�n����Fb�m��3�#��>�S/{:��D��(|�\��٦�2�Bi�݋�3@G�M��-O(�QBP[���&,�!�����כ�Qruʠ�*L��DH_��w!rY���<�(�;ԥt���<
����(��,o ��ك5�"�̬AO��_���(agtbTX�W�n#��P�$ =��Ł1��iwlu|ш��T���8G\(.�eۂ�M�F�'jL��pg2�$�ޑ���]��y*�����%��fi�_G���:�� ��Z �Ո���V�M��ƛ�i�X���[w����V�����~, 8@��TU)980�����)5��b��-x�����z�Ѱ��ƅ�-�4x����Qn�g���P�[l�-���IB����J�3G��'��H[�#���5/"]"�f���K�|
�����֕��k��gyq���� �rrr��������6�L�%Jn<�{@+Z�����B�̃�G�±�a��^y�6�#M.~%��w�� &�U��K�C�����Zo����ݝz�>,߆��O��ٺ�ϸ8��z"���h�S��[�:ZP :T�a�X�Xǈ����{�̮�vD���_����O��J�)�@P"x�,��,&��s��կ�2a7a�����;��٠�{������$DDtb��15�ޡ� �"��T�р�g.x2��V���B>" �
2u���aœ��(V.l�Z>��I��.*� z�ɕ��x� :a�E_������@��@Q�_�̻5��?�����K�Go%��-,�D���55����]s�H��E�K��kV�P`�s��]�w4)NҺ���1�`�odC���Nʆ+KR�k!��8����~����'Z�b��$�K�]�K����=���0�� �WQ	,,,��1�  Rna���:�`,���_�z� �7�o�ZvA� 8�qV�n9
�B��zov��qd���t��8�Ҫ�yBM�8�e����#�� =��6efvf�*�b<DEE��V����k��3j����u�x��z.���UF~!��1�����>Q���PL��_���)���,�Mg���4o�f67�.--��RKHH,��`%h����Ӈ��w�� �մ q�:`�1�38�S,�A��a�S����6�>q�Fz#���+V?y��������ch1����M�aI�1Ѻ�$�r楄$������\Y�:S��@�x�|�f��ؘ_J
1���a�z������:��$��W�b3���/[�X�P1�d0A%0"�`&\�|aM�h��pܜ�/&$�)��*��N(@-����1��L%gL�����ۆL�~�y�_������f#fR���K@�5��}��Tܾ*�|+�*�ؐ��_��k.�����h�w�M�CeI�XA�R>�y�L5�B�}(V/�x�7#�S�w[C<d���;*�v2qo��X���z��y\��_��;���w�
�K�j6\�l�6l�sE��5;�r��m������ѡ8H�k�M+_�r���F��1�E	��~�H�C.Kr-gZ�&��mD��ba�Y?�� �I�v����z_�\i&�.[������?�si*�v�J������ʇ�`�ep]�}^��"P��΍�(���췐qUU\TC{vQQ����MT����ߊt�qq��k�����M�K~6�N-�����r!��I�X@�Az�x	���f�Z}���F�d��������K cB .��1�!�
�^��u'��� >_����ٽ���j��:$2R��K�ׯ_�"� ����y��E��- �Ի���r{�9RtG0�S��7Q��<N���j�[�D�c����-�ݱpV4�����z��>�M�YW>NvdQ�Đ������=�~��+����p�[/M6�r�5D>T��������4�>1�nz:D�Q*�l~]�H��a)V8��5��?�F�ð��iZ�d�&��ʋE�o�^9��ޙ{���<B@ߤ���1�.5U����%���
|V�U�2r�7ic&�DA�L0��AW�fmsQ>��Y�{�[*ib�͋��җ4�����mG5ď��*�O�����!/.�<��`�ջ(8�=��'�N���\3U��r���b[3dh@'a�}����rM�Uϧ;z=��v��V���W��[����������&�|-������cOa�_Z\ol2��ʴqq�N^^R�g�����k�o˾�ON��KL*~B��b��4���hCW�l%��D�b1�&�1����U�YSӡ��l�3z�M�ndH�<r9� �3�@������&�繁T��q.� �ST�B#�r��_�:i0�+�O���6[xy8�B��`���6��Y��6��@-qϜ��ÏvvN�tO]�i��$=z���4��y
ܺy�3Ɵ:7<�O�>�4����P���V�h��;|�DǢ�a\����Q�r��D�+��=�� B�Vk=�(�w����
.)�"^+l��d,�>��~6A+@]ʰ�i��l�Ooޑ$Tv��{��V����ƶ�2����]�Q%s�%�_�1�|������S��Q;�A�3�V��. �;�y�#�"���ϴ��"-
��jK:;g�ι��-ȽǱ_�p݉��u�t��de�܇�KşqppB��_��_to"�I����U446����gR/k�m��d	a��o�Y��z5���ύ]�z�/x79f&�gx]� ����-������W+�
������-"슾^�#tO'��a�h�S^��R!M���|>ύC=������]� ��*�+LF��1׹g�۶����G�0�_�(NŲiZ��^�Þ��̛��"U�ߣ�U@�N����a��u�#_�j�k�lS��N�G�����G���4J���|43����E����L��6�'	�&1�<�1�B�ׁΦ�{���v�(����FW����r��t�)�k�@���f��C!���xH�=�#�;2��]y�)�!�/����FQ�LK�-�Ϊ��QX���4��]JH�5�71��^l�o�ۼ�A���_E�_?�m��,��}a��`��M�#]���Y9�V�G�FT��x��ͼh#�F�6/�D�c�M��co���[*�WB��b�ۡ��E|!���gF�iֶt����IR�{��P��X͹�=5g����P�1۵QG9�����i`�/���4���܈oC��J�2_�d}���B��rN̈́�s���w�=���Wp9G��q m�@r?
r 'V9�����a&Xa���đ@IA�D�������1��E���
0�����@	���qt,�ۆd�돾�.����}z�(Ճ��WK�i��C�݌���:������>���ⓢ~��;��ëO�O�l�&z�A�g�{�,�UH�&	�t�v�ѻ��355����$''+��F��������ܬ�H���	AH�����D���%0Rh�0\f�ȉd����g|&*���p/���~�gŪ��I�Y��~eݓ�B�{R�<ժ����\�����7{��A�k�9���L����0�j�m���|`�gd�ۿ�$�R۝|$����ˌ�Wr^0���Ld���=�4�I]�u���b�޷c4��&�ƫΏz��)�b'���;�}u��S�i~NW/�<��+}�I�4k����ޫ�.i������7�%瑂���3ǎϖ��4=S�&H���7��ս���U�B�ֻ6nMǷxd#�i��cj�`�0���GdjIG�Ô�����F�Xz:Բ�v�up(S�������j�&��kj��DR_���e���R�|�p�:�X�ol\�仠m��Q�5�G��~�@�Y���j��6���+F��-j�� #[��L���o���dd~/��'��;"5j���	
@2ED\��QET-�侕o����?9ۈf�\}Ƙ_�6�>q��CN�ʵZh=`������7mǾ=`d
��ӭ���QT���]��gt�E����=}�ِ988���Y�������P�t�%% �*Pk NA{�>s�A��gE6�j@���yj��U�j��ΐ�����1j6%ػ��Y�+;WL[��J�[�Sgɻ��V$#���a��Y�~l���+��f<��0��P�l�Y���7{˝��� ��ʈA٩�:Z��NeD��c˯6�:v���Q�f�1Fp6v;�4/F�?`�.$w��*���H]Qʻ~9�!$�Ci��Ұoê�O'�p;��q�A>�]e�	�u���\����5���!WyC�L2~ep��(�+9i�4\���@�F�<�'�X�ԡ-��~_^6?%�Η��F�w\�c���j+]ٹ �u�ۙۃ��.\זq@�pF\9��r}���h˂Z��j0�w$o�DIɔ(�$Ȯ4`�=mE�Nn<�#�PXU�@��v�v4I��J��y8��I����/F��aw�af�/*穧�˳=ϴ`y�����QE�TT��~��~$1�.Jv�=� ���i�oA!%��`m%�܌C�t�i'�Y���Q'4�v��fb]�����׌E�_�փ�ż鵎�;�l3O�|���䝗�^������~��� �n�a��*޾�f�Q�l֭PS-M���E��f,�eN�9U8׆�q�*�{w�H^FQ���͞����^?�`�R��YU� L�</���p��>i�:��b����4�%�/1� �P[U� �dA8'�/.,����wUuV��0�L��������'z8��3���Y��g����{��넍+���FM�^'���S>�EEFv�O��wq�j,���z������R�>>^�37ۜ.B�<��F�]�*�<��a�4��q���5K!���+񒗽O�"��ƈuuٞڲ�����F���AAؕO�Q���ݭ{6���'6���u#=���t��5j�7=����zm{���y����0w�\�3k�]����s`�}*�I+���:�#����"8��s%íƹ�yl�e��TV@�8�?��)u���w�aɶ�6.>�����ԫ����5}�Z/R h�-��t�O�4B3C�l|~O�]����Y�]?�aqܛs�� �8R#G�-�g
M�	qvMC�o�Бܵ5�{�V��*w�s�`]���v�w]^��Y�#u�La2��I�.���<<�NNN�VVUw�ZZD@��W��g+�sprb^'6��y� �3�i�l�]�j�a��ˊ�7-�V�.��V�s7�����X���>xöՕ\�du�G��ZG	0�\@Q�� �;8�Hod����9��u�LB�0�o�����by��I�4W�RcB�|���=���յ:��7�.��ɭ��jK�0��9N��y��d�Z��;vh�n��> ��2�������4�_k��I������\;�j%�ļd80�g�����4ހ�To��wn����꬜��������d�m6�mꨴ�TA�=�4a�zŲ��߿�*���=�l�___/5�ʷ��E��\z?P<""�u8��Xޕǳ����V�\�:L��eh���z��(����{�7�y������>�-��@�OOcss{���1����0S�7��DǞ`�S	������}T�}��U�E�7ׄ��t�T�����K���/���F�zߠ̎L���2�3F��T�쮗\�Z
�xo��j��n)��fO����@�}хyt���ʒ��%'79��i3 �K��C�ndBX�<߮��V�L���>+3�ku��-gqg�*3n�\�6LH;�������c�+[$��0.���"|"U��ݡ4�}���ň�j�Xd���y�����R���������pzxX��*T6������ϟ��]٩v��0�t��3i2ʽE62%��c_|�p�3���g��O.B���+!6��P�!��搐ݯ�\ �#��#j}}}�|����������!�M��+/���~�]�-vVJ��Ò�\X�r���eߟ'�Jfj$6�`���$�U6du�`dBf�A���О-1�m��񿼙M3{\�jCBK�?.L�*	�N �����)i�������$
Z��0t�~�}#P�@�	8����"����Zi�t�u��W�h�,z}��p�{g��H��	?�{ 䵢�6\��;\�mԤ%!�bQDv`CcK6�m
K|31a#���'�5X����?o����3��ޡwf��a3;'��H��9�d���pe�Y��'J�mn�7kcJmI��r��{����F/�&��&�τ���Z|�0ZjO2F�/�0�x� �0�./y��P{��~qa�4G3�XG����ͫ�#��t@���út��2�"T�M�"?�ћ_Ω��7&)����o����xdb	���=�`���C`�nC��i�.5��7��[�^]7���
�A{�+��������s�J'��L�M��(/~���4�*#�&�c]B;EІ�
VS@�ַ��w�A�g�>�����qG�K��S�"D'�oHW'4#Ŵ��GI>������Jamʆ
j_����bu�UC{Ƅ�$'/?6��IU��:vu{1��Ϫ���R|�� �8��ے��<�5@�Ƌ6?���H.��Bv�V��XDW�nU�09k?���Gȼv��G��L~��BL�BV�D�'�ɠ�f�(�&��jkDm,$�t���ۑ1Lb�\;w]�`���ǽ��ZbTOjϐ[��pGǛ�u?���w��R
>�<H�J�aU��V_��)�#d��'"o=Q�4n�]G	���z\I W�G��M��z\������u5�D������������p6�-r$�!nH�)4�ڑ0�&����A���=�/>�J�)ֺ��ՎҴ�K�6G��mE�t�-'+o�����o�GOO�NN�|��NQGn3	�~���*0z��^8S�	��/��0BѧW��&��E@f�rU��p[�Z<\��dXXd��g�����O�R^g*�FȘ6?�7\�I�!���#��̄��E��D�7j��	�<���e�v���#�H��}��AF��|�V_�i��H�����~�'a�m�����MC���Z;��DbӚգ_ҧX�DP�\yt������i���$��υ��ѭc�D�Ig�٪��3OXEj-�O���MbDP��^�Sͨkm!���&I�?����(u�4�L	���r5Ǻ�F��t�����]�
,�&R�T��a�S��!c�FW###�XX7f>���B} ��L��v0O'/P Ú��㣅T����o�6����(k�46��*;tL�f	���Ro_�]z
3t(�I���i������z����p�O�M�P�=�L�p�Wv���	lE�������`q�@�r̎RB�*�c���h?�MdTkZ��w}N�q��eYcC��
	ڍ�q̯b�4jy��٢*Am�^a�����{@-�Y���t����Ň��պ��z�b"�q�'EM�|7�G;!�C��(���ظ�ڭn���d�@q��g��`1�E��5��;M9��u��F,�+d����}�]����6T:@�����d�.$K	��	��v�ĉ�oZ�S�UUSCEKO�K�o�zE�K���n��V"�K����n���ɷXy���$!�n�"w0_�=קR�h�;	���LQS��ľ!!�.��7���n�3�y�)�u�N�ϊu˃	9���UGũ�M�C�p���t�^��j�j���B�^QqY)S�A]���rؖzR���K>�n<�x:m��>��=N���]ϸ��L~g� _�PK��!�;�T:�		���W��! jA�U��ޯ�"yᦔX����L�����A��|d�?�Z�j�k�H��x��t$u��botRW"�D���5�r���� �s*��6|LЂ�dBVj����G5���t>�\�P�Z���&$�w�H"�h��{��n�J�s�jۊ���	�Rd ��
?���"TRW��Ϸ;�-Rͪ���fc>J%-*?A���x�N�9��l�CN�N������CCA�}2璌�7���V������%��%��=��'���)h�)�E����)*gO%l"�	S`<�����w�Qz�.{ø�f�`ְ�	��R�C;���^}���DGrc�Ťx�+4^��9�����@�3�B:7�Lқ۸������r	q�����UT�I�"
��!��J'\��7�����a�n������g�pb�QK �]�zx���Y���\.���I�z�G/:{ӻ1[ a�S�De�Gم���R�rr�����!!�/��R����Чib��~���)%%�:33�����y�.�M�骶>�k��p��޽l��!62����Sc��;55EGGg[��ݻw�a���|_zQN�e�,������'*�y?��1R�s��XAp1W����J,�� i��La��k���Բ7W]���S�H��,]��v�yT�����MO~���B�443���%w�W0i�mƓ�D���DE�5ײnw���ƹ�]3�5�O��s�{��	M�����\�>�4�5�^�{8�mrb�О���tI�4
/Fs��Q&z���|�=��M+r%T)�kX�`"��:�W�Q���ƍ�o�|��zHO���?C�|�.<�.5?��7����ࠂ���je*�:n,��ի-	��j���.b�j*zЉ�SJ<_ҞJ��$[�8�����ꉨO�1AE���W��D5��X�&'U�E�&BCCMMMK�� ������p��]��4cL��uV�*�W}k9~08}�mq��1zGs��ݳ�j��j�ԒL����ݧKt~�O�5��be
e�+�Q��j;آ�b	3Z��V��;@�1 e2���tdcgl��:��( ��V��v�^��@Y�r$Ɵ�#�L�$2PK����!�O"t_�M#$�,�6����5��L�`b��مaX�Z��Npl�N�q� �?�a���냌�ʪ;3�P��yܜ��kW�G5uu�v��O�2C*+���{{�MNO���s�P��̑O@'#;9�%��K
RM���Y B=fV:�O����0�r����Ӏ�^���ƴA�b ��#��f/��ĵ���E�D�����G|jt��M�UC�� >bT�0Ht0\�S�*�Ԏ�6��߼�#81��Ba�N��*֦A�e����ȜU�����v#��%�����`X�&��Q7��i�k����"\��5Ta�pzU!�?e��`���wx�Y�{���!U��ij�i&#�}�{!�A!(�b̚�o68�y�("m����Ƥ@C�[UF�^���U������(㬌����a=Қy8΃��k��`��g�ʝ
5�Hx�sS��je]:�\�����|g�}�Ud�Q E���tg�������٩���A�t��Yii�]'{�9��߿�PF�9�[��13o�l��`�t�C�����DW`�zٞ[L���F�.ք�����	nbt>,m���[=]��p`���6����A����MQ+���M��������h��(`K���Kg�@��]}Ӥm��� ɤϚ;ʤ��,��N�k3�wl��*\*T�����d���[������<^>hw�`t����2a�ԎV5J��tl(���&S�+	Q�����̠�F|�.Y��2��)��Z����j	��d$�+�r�j�Tz롌E�������Ζ�����4���7;TH*�G��f��8�ML&f?�H�]F��K�)N&ڡU�9��kjuI/��xyBN[���}fN���=9iQ���`r���/�Å����)}�P��`�=�lR����>�
-wwwIh?�;�������DB�#>n����@C�O���RK�Nl����"%��_j��
t��|��>Y9/���R����fh�� �&##㑪��t���8%?��s��w�z��:1�����8e���[�u�ɴՠ�� nX�ޝ�62#F����`���K���59%d�d3CI�M_Ug��`gj��)�Ľ�O�+��;��e��!�籭�eU��_��'���-�Yc��̛)��!���|V�Mꪼ��y�c�tBN3P!��#���=
'��WR��^��Vc�*(p�x73��xEuBvW�n�w$�|�0�u��wu�����Y�>��!�^(SF
r5-	�9��^iAq��+J��hv֗��pN�y�vU�8�h�|�c�>d��H�)l�a�90M&�m,K6&6: ��ёK�D'�������#�Y��[WG�䔶g{:ě��~��
�l1C�Y��vҌ�c���z59�Y�jjg��'���S������h&3:!1�=����ǜD�T�3�"e�iU����xio��	�E˻U�/��7�ذ�������2�����Һ��@_.�
���Mx��D������×��z��'�2�8ne��r|y���&u��ۣ��k��oO[�O��P(�D�Х�L����ȳ3U'��}��\�*#��v�7�,���k�i�pӽ�˜���p
�LX�벏���/O�o ��7R!�����vf�F�mf��&_Y秵��w!ȝW7��Yۨj�;�8�ý�*a`q�gts�;�+8=���n����ں����G:n���ww�\��C�gQ��5�L�5CF}�.�列k��,���$AROG����[����P��a7��f+��N3���0-_e}&$:x���b%�O,�y"sG[�3��������2W��H7�$8���x�_^�4^^5U������=���-F�/���o��쩎�⪣@��U��N�1��Z������jxQ\P+�P۵���\�(����M	�������J_�]�6]�������?��2,�`���wNp�����B �{p'@pww�K���ݝ��fs�}����23��U�Ω��aA�����X�����vf�}�VoSxu��q����Ep��9���+�s��*C�^��I�?��{���Ũhg��gb�]��]�&�Aw��:�Q
��tX�߉ M�j���{w*G����>}|���h�����?t��yM7f$苿II5�	�#qT� � �����gQD���X���ۭ�Q�-[9� Gm$����HP�j�&��ܒӢ�׻q���\h�1��Wg���'T�_|�~�]��}����(,�*�>�-��҆���:Y5d�(�x5��T�Ȗ��K��i�sӞ��J/b� ��>�Po?�d-�
k��Ftը�#�0+�UW��^ ��b�� ����9C� u�M��~v(�qѯr�b'@r �#-��>dtx?�-�I�Dl�.�`&�ѳ���4?��:]�a�>�0l4BhBE�Z�ּb}��u
��o�ZY��0��0i�����J�^tr�e�`o����`�������;��eg)oa��|j�k]U�_�\�l!�����B��R�rA[[&8����:���EE�{v4�_�`���_�Q�)�X}�o�X�A�n
E�-��_�f����W肳��;���v�-�T>{���F��?Z�`Vݤ޴e�4���?���F<��,�d��<3M�ꒄ��.f�0Z�.�f���;"�a�GS�GS��!v
�HՕ��խl�}�W��XE�ܗ�呷�$*��/ZO��>3��6�U�F�4�*�XC����Ҏ=�����r�ۼ>����w���Z��8E�ԓ��~1��yT"��#a�(���%�q�3RA�υ��VT7;��2�a��P�Ͽ�x�i���Sd��0�"��Y�����]�HG��z?�F���/����r�+_�AOk��,���%����@�b����@����ͩv���m<hg��i3
j"J�h��h>K݃��"�O�V���M�4���D�Ϲ�i�W�1��򊉏����歧z����z���NYW7 ��L�f�`\�����(����k'
���C@χ�l�։�b���4����a���H���mx�h6���>��M�p?3���E����BVĩ)��h�9���K�JH�0W
��n�h����9�&4A���Q���6:
��w�Ú��`k��0���\��o�Ff7�z�o�9R�ng�E�z���WU��X*��F��~���s��:Kc5q�w�r�?|tS�����,і�����������J��#NiZ�In���<8��	<���.5���kdz=�,���z�_�އsJ�w7�qdL���;�O����]>P���J���M�f�8��]�Q�=��dB�y�}xh��3�,xE��޾�H]]][O��5��ht�(ʴ���$�cWda�-��0�T��[x�=w�0q� �[L4w~ס��~���6T��
�Fa�x~l�f�����U������s�WW��"qv�*`JwOK�m�:-��5���O�ѝ���zU��GP!���2��(x�ܰ}����Z)����Fv��z\� ���@��ɹ��ef�u6���!K#s�n*y5�ԙ�ӷh!Q>y�|��G0c�z�G�S����{G����C�k��_��<�KI��bNN܌ⓟK+��h�oκ��s��/�/�O(}�G�Y}�/G}�V��Jm>?��&2�O�c�[}UP�b�Č����(��Ox}����Δiɥ�|SJ�Ob�.�Fs771}U)���st��Ӭ.�@
E ���/m��_ȗ���v�x�.O�;
D�QoJ/��Bs�x�1|�Td��h3A�q��n93Q���f�����\�n�i=�������$��X�$Қ��ɀ�Rd.|���L��ƚ�9�P^Q��U@�Hx)����Hp��n����]�^�M�iC�!��wۮ��{������ȋO�>����
#�7�������>���o���yv~?v��o]�������++��m4��{xȻ�h)�bA	�ͷirn�'��)%l^�։�B��-���D�T8����h�o���ͯ�Y�W �خ� �k;�eO���<f��0ܤ��q�Ȯ���ӹ�kü��r��1!]����+��µ� 7e�R��B$h����f�!~CSdvy(./7=Yjz��9������ù�u��2�$���9,r�Y�'���74���$� ���+�R�8�^\/�ʣx,2�ٙ�͑j�I�˭�I�"g<����L+
SVq��u����N�+󣛕D��3��D���]�K���ɤ��P2t�Ņ�f����*6F��o�&!'��b�I9iqL�u4��:�E����R�=!�4�;-jϦK��7�V��_O���:OqC������#R@� l�A뾯<��@0�����B�����B����D4����B��F��&XA,�(�ӻ�`�2��!|b�#��mi611�`���DU���$B��@���������P���>�k�����U�S�'�b�b��^�o��ŗ6�X�;zH��>
Τ�^l�F��r�������Y�U;��dݟ;N���ƤUC�΍F���t�_Nl7�p?��Q��{���vI`1��N���w:���[P�?�Ώ����K����jo58������� x+���G���0�t�tFjBCɽH_��J!���	��ءG�c��qfD;A_�~��T�A�v�����������p����c��+�����ss㷡�Ө<H�1���Zy����Y�� ���u��u�y�M"#t���y۰,I��W��T�iV�͝c7�6��x���v@�
b\%����Nw�26�{�;�P��Ȣ�3�ғ&��Gk!��֏r�i���mcӍ����S�C4��DU2�$�v��9l�>�&�H�^���6~�.�e겚Hb�yq�E�m�ᡧ��EIؠa�fX��:�r�"�c�CE�Z�Hn�9s�a�'x���������t�юD`�ҙ�rv0����K�lӥ]0:�w��Xs���BE!�&ȶ %y�����FS�K�W6��Ӑ����g�Ozz���8ݎ�b�<g76����6,�l=A�z� -Ih?|7��>p5Iv�(~�q.t*n�:k�gP<�j�k�5`k5�1��a�n^��h�d��<!=�G��	�����ٚ�`�t�""&w� ���=8Wml'�"�o[��9J]=J��� �d!$���#��s}�Ɔ3K;��Gw==��y�����E����|]����)z���LMbn�$2X\\�D��p,��ɩ��8�8��~bRЖ*Zbtk0��ލܵ>�#�I��k���%����~{�y��Z|���=i����$�qk�:(���*?�W;�����A��1U3�����zp~~
�h�Ux�ӗ��$'ϒ�5.�{"m���W�H&��.!	k����QW�
��:mQ��?b�r:�X��������"���u����t �5߾]�L16��;Re�+��]��?�� ww����%%���;�mZc������Y3��v���E���\-�Y[1.Nb�P�X�f��NZ��3~�V��߰�h1���ҟ.��Q����C8��ra`p�,1,y�R_Q�vӷ�zv k�� ��*M\��Kn�{`Dww���i�8a"��(�)+cb�)�'M]\�@�B!.�D�GB�kM?�w>��9dn�2/�,^��h�Mf_6���N�h��]�b�|�v�ݞҎ�h���P2'6Y�8��|M � WE3C��}v}TZ&�wn˲2�����/���.'�^�jj���r�'N�v>�\L`=gy���4�����r�ߝ#P�p�ͨ�%�c5`�k��g���<�
 �p>�h|��������`���$����{��@�����.�ʌdk�[*<��|��
]"F�Ʀku|f�d7ؤa3[���һ����o�'�SW�E�ԕ�@'�!��oC�%�X�V������4$P�"QnF�}I�!isT\�+E��Ú#���{���˗���1��s6�#A�	��������k���U�%W㐥�N��{O���kJ27��d��н��i ~ن���K)[��R�D�/��cy�$���l��!�$�(>�ef$�zY7����z��=K�P;��?30:pr<+q�̠Pg�R[G�e��vY=Ϋ�i�]5f�l���ݱ]q�&�y�=u�࢙�����1]R\���@1B�r�l:��yꡰ����;�"N,MJI�}�xq�A1P�S-<�!s��WgaW�.��/��5ڰ�����D�Y�O���[��V��b�p�T���}�y�P(8�����E��w���eCjj:�lV+���Y��g9"�?�3 �ŝ�K�<$�g>Eͣւ����+h%������ɂ�N.߻
1DF"�8[x^ń޻s�>��;���h�v~8I��Y�d�~� "{כW�/m��d�v�p����p5���	�����՞�]PJ5��պ�Ul�%�駦�j>�+��D=2_D1��I��0'�ߨ'��pS���7�i-����i�O������ش=�7�!�8Χ3sM�=3�D�<��-��˵Aġ��1J��JS�[w}F
0��x�9Pq<W�h�d�}��ܥ)"N�UziX�հ�m,�(�Ti7�9.n���-�}y��)��3+z�NFJ�FMju�| �6K �Xԛ=Q�p��>������Ǡ�k�b�/�Z�-U��*Gs�eO��H�6��d�)�6c_��V�;J?��1����M�aFOԻ7��}�y�#�ȋ�؝s�B7~ரg���!YX``t���`4��a�-Ш�O������11U��Q�*f`	&L��'���ffl��JFu�0��&�E'F�%���g\L����0�1��x���6��et[�$�^\�Jp��I���9ܳ9!+����k�}DP�����~����4���ō����@���e��a��Jf�W���!��|Yz�re�2��?z�����*�۞T]�&2c���F�q�w=#G�����*P}��ŋ�j}���ǂA��5 �"������5K�������P; 儯�M]�k��Db�}�yާ[VXb!��9�^��x��NX/�Y��$0kן-�z���o�
 J�h�HY+my,��AQ���rb�tM"완@�VW�F�중`�>� �K�f�4���h�FcGo1B�~v��D�4�a��VT���y������yv��!�ijj**y�� �<hUt<�{?,��sϞ]f���ڴ'��yDB�FPTDd�	74d�c��(�GW���:Klѐ��4�\��ղ[/�=_���A�F۬d1�w�Y
I���ͧ���C׻�Ħ�m��ݻ��n��t)���m7D�9Fo��G��h��Ա��~�ߺf��/$��OT�P���󤾕P�sJ_�n��p#�ըa�V�;���������������ښ� ��t�90�%�? C����k���7��Ip���z�b]��gl��-6؀�L��'u9�Y����P�4l�gimm��B���oX��3Q�����G���y�9��ֆ��؉�~�����>l�O���Q�����d�Y�}E�����I�����*���a����K�V���B���J���v��u�vӐ�mu��NK:���~EK��BP�MSx�H!��nlaA��GX�ݑ�����9��B$9K]]o�������7��g��L��i��++��HA���ˢ��q:���l2�@�0��~����0� ���������g�.,,���|{D�t�׬��Np^J
�b�ҡC	�
EO�o��?��l��~��v<��3���X��g�Se�+v�y�1�����Y3��޼�P�z!=Z�@!]��`�)cc(�ޠ6	���[��|��A55
 ��C�8��"������'8�0��i>#�;��X��鯽�gk����0՚O�6��:��s�s��_\^j5�R(��o֚m��'̈�0��Gs��kƏ��f"� G��;�Y��sY[ox�+>�5nC�-��r
!� ևl~Qu���lxX�$	jk�����勨8�q�V[.�iؾ�I�nx4�i��\'p�q�����
��/��M��jM&:�i�a����	�b��LȂ����)� ���&g�q��o���#XLO2��J�~�gx�5p�皋���cz,����F#8c�v�'���-�?��SA6�+����%��4U4��q���"��3P����[@s�  ���|$h�O��m~s��t�7��UQ�6;�^6V�h�R�^޵{i�&B�g��c�+r�ε��!u��8i��N�ˎ7��f�TR��Y��܈��"��њ3q�=�Ha���v��h�Y�!QfEB��%@�����j�L~P�Y%%2�� ̈́��������v�C�zu��/�jqfN�uN^Z��� ���7Ǆ�O�v���]:�ORQ�91���O͢�q�j�`�4e Cl4�z��ui��8�T283Ƽ�өf��u��f�0\܀�����]/�ò�ۇ��	c��s��f��/�˲�q��b��J4[�h"���]g���P��^��wN�'彛ND!�e�̑"vj�쇾��<��ȃ��:����'ϫq)@�E~x�����7͡�FQ��W�x�T��m�`#�ŀRg:���?v:�]©m]@�*�1Ɗ�M��$���g)�<5"j����NL6_wU0��~k�(�W��L�V���"�fh���{�;��C���e���|�j���:���e&��������6&��,9)\�h�Y-4�՚�MQۦψ
!i��F:Z-���$���������Q����_�-w����***�M���~r�4ȪO�|-l$6�0
���cLd==�]i�Ъ�"F#�{6�A�����1Ә�$�4����ը��'|22��|��м?�8:����p���"�]g�Su�ZP�!	Zn	�n���M�ݎt? rC9�s6�	f�um@t���\ݧy=�(��'d"QH"˫���ъ�0�:꾺��C�D�!���k�����gM��w�b�Z9�>O�eZ�𕳋�f߮���R�B_G_z6�M��A��	o��K-)��3l}��b�O\3R~��N�9�&[5�{�Oc�U;"N#��6ev<̻�SoE�J�)����a���V>E��iD�Ю'���)!=����u���}������I��G���}��o�3�/d?z��y�wYq�����A���yX^a������V��P�s⊢����a�b�@^7�n�ˑ��8tC�������Z1FYt����p��O���u�6�o�.���~rF�n���*
Ž��o�6���A��C��~� �y-�K�x�M�m�H�XźdaP暍��j�\C�����]��6��P�N;2�J����	�-��0Pe:E)�W�
Fڶ���Xe�/ �2�qFi�#C;��Qt��B9�n!�z�/��NLL���횥�h�/Y��Θ�&����_���e_~1�s∢���BK�+^"� ��q�S�>cz�0�;7*�a�a��?����jʫ�p*$]��P�3�rm�W����q�(���H�sN�����J��hux8j��ȓ�f�:��j�{?����5(��MbDmEQ?���55��q??�f:3)���j7Xo�ʲ�k�˿eT/3 �+����j�������-����Xag<���\��R?M��@x�xh��Y�X���8���8p�rc�<�}Z���]��e�7�0B����f-I��j
%��e�{��u��rގ�0�����׀:�ݸ>�A�Q6 ���b����ߔ�@����9Kj�+y���)y��`�;6�*�e_OV\��X��JAO���`��V+_�d�c��b}��)����.ß^)#ڕ�<n�{y�49���)&�z��D��ؒ�n�E�zQ��g
O��+!Ж���&�سV���x�z����O❻*!�5�������%�IgV�e���]k������7�'�����^n�-ZVl[�V�����Z[_*�j	�TU{n4ĸxJ�^ZW_V�ڽ�����:�T�EM"z��kRٓ��Q�P}�2�D������i��� /��a��y���n��x����{�A�H@W-^-,m?�!ˉ�����+������Kx�¸"�a��/��z:����ۉ�������ҡ#�X��h��㑹�VP�g2�T��G��|IJH>k�Ո���m�?�Ϻh{��G羊����E���h��^l��>��d��0�PUN2t=t�e[)�RK�p�L5�C���7���wsX��Lh�WLʪ5���js�(X�-5��i�k��,�B+�.���M`�Ǔ�M�K����5d�#���z#���[ 8�ׅ?9��9��K\�k�鳻Nኯ�&�CrU���@R������C}�Y���:����p#��O�O��Z�zW�d�(l��J��h4��ʨ ;~'���i6ѐoz�D��P#��Y��a�֧�1�� K����h��Sw�9W�n>I��3�Ǣy7�'�T���*Ջ�s��.z�a��p~b��г������u餳��v�ɐ�C��{m����_����������Q�a�&�>�� 1F�ޛ�����.'����-S�1�^kRN�?GT�o�D�ƭXD�'6*Z�T��"I�[��IUq�<q?�xf��{�o�2�?���GB��L=�{����)�St��.|-��MNoe|�a�Y�Ԕ��Rj"�ǎD�W��	�����X�ho������4����ag�U	@H鉨-B���ϓ\��+5�b�s۪���++c⅛*�?T�nl��/yT�U0Y{\){V�������_i�,D�{�͗�
���{��t�@z$��1�EB��5���e.$xގ�ߝ���cl<�A<��H�8уe(�p� u��smC���bW�O\S��3�:�~�]��e����J�E��I堄s;�Z�2��J@/�[��Zu!o)�3\͑�] 6����? ���0�ف���T��lLK�u��a��"-�ݎ9p��[8�6@'�x�x�;zz����w���Gz���E�"�d����	8T%(f-��Z�w��:�0Hw���f�=����������H������ia�M{x��L����*:*ߣ\��)��u{��q��m1�S��	����dǋ�Z�����ʤQ��q��++h�	����0u�B0+/������w�	̇��Ƶ�I�`����M;�Z�<�U��g<����BXވ���/�$@m�;m���&&���ZS̾�_v7Ƥ���U�z�`�Ʊ�ͥN9ç��a����->>~����ZBy�x��v�t�J���J�WeO�a6�sW(B�|E_�0$�#�?u��/O2օdY���BB�6��y�6ϣF�f:���ڰ���������I�l~�]��).\H�Mh�zM�MIΏ�*��2�ɩx��5�Z��w�
���K�o_��
�8BB�D������:�=+�Y[��F�)Z����&������:�W4Rv�p����}:�Zi�3^�Ck����7�N�U��O]�CgǓv�z=���	��
�=�=���eKE�E�m �wPX2��շ�zL�`l2r&88�R͚��'h��ά6������筿dt�LԻjW3N=���XO:7�v� ���� 2�H�W��(�<��"����Ug���&�]��E�Z�Y!-��6 �_�Vј(�]�g�B~����	|@W�xm��ҧ��p,n\I4��#��2Yi��!޹?�~�JS�~!]�U+��t0�3�K�/_�@���f#B�����s�Gظ=iU��1�4;���5��_]W2q���O-�\�R~����(�҂z춗��Q�t"�<�ɼ6z]����%%�T(�K,�l+���͈}��i�<!�r˵�ҩ�q>��E��{��u�I��7ԤY��Vޏ�����2
]1JJf��-'�� ˳.��*�7����*)lj)J̒���F;������T���睯�8y�� ���2CKPu#-q�(��82f����og�"�k�7�¤��$�}�'+33}�BB�tG�ݴ3�X���ts��"�<q�e_��On�!�y�H����<I����T��H���"�B��4�ϥt�kv��\��T��1D��^ŧ=TU�t�+��TYQAKD�T����-}>=(��X��wXvJ������]HE@�ijoɟ���,���SͶE~��+2 ���'1�?2_��o��������C-I����[���2We��ׯ_Ir�����˽���B��Ă	^�&�t�h�
��¾L�}��֐iX�r�A"xcp��,>��� ���M�q�iW��c�]����A�D^�.��XO�}��yw��##@�B���Q�K�2�w������ca��5D���p=�� i�Q����Yw�h��	�d\��l+�dY��b`̡[�ʔ�����b�V@@��<�Ô����\>WJ�u�\E����0��&�y` �:��Pw�Z霮z_��w��>!g<���i�y�j��w%�ȍ�ӂ��ųrm��6H7W��=B�rnU�Z�,�����&�QQ.?�gX���v�͓��S��g�Z��לn�"�͍6�I��cq����&׋I���-�>1M9l͍�{~���9gf��~�7n H[�v:�Q)�)&lY�4�ೣ���Fz����R���=ߜ���������r-o����l��X��=�_$���6�����v3y�ͩ��]���t�e��m֏j�m7_�+��!�o�ȟ�<���<l/Xv�����cA���b2Y "�E�/)a`i���K���ϝ����d85MDC��RM��Xõ��%Tp��#�|$�G"�ݹę�z�F��v����|���6)%����֦5��>,՘��JFv���{�ަ��1	(���!3�Y=��8Ō��jE"n�/��il�u�#�*r-�1�<�U<G?��^3��F�p��ʜ4!̊<������T�#��;��~"�XŁk��e�1���RPV���L���Xe9[�����A���ȃF&��&9kWS�A����p��-3t��K�p�oҌ�h��^��Y�׈~� !���n�����m1��A"sך�Fb6����غmR�vCM�����s>A�#h�G������N�vP�/R <��#ka]f�Ps��y�Dv
q�]�8Uv��N
��q���wCFV�eq̌v�d�^��ʦ���\�3�;@�%�����J���u��
��� �n�T㿈7W�ڬ
A)fT����>�K�޻��Ђ�㹎bx�hl���o΄-���o�7�d�S&Z*4P ��&�M�KXy�)6m)�^���}��M�꺺�����"�}���i�c�SY���`����2O+�?���Xf��jG'��j���x����B7��L�>�x��w�-�6�����ca~o�+��IhkkO8ض,�LLTQR��؜����Xu���|�%������s��t�b���MZw~�@�0~#�/�*�*js�^��= ����}�N�1:]$�*n]щ�>���IM����)�]ϻjjj��4Ž�uV#�v�,pI0`����G�'nbO���̦�,��⑹���W��	K�٬�9
�D�+}����W< �_�@D��n �`�W)�i����'췣���Ք+�lF��E��
�R}o�F�y���>��C�%w/nJ�N�����\�dF���h�P��'ł�H֔��t����d-�;� �Q�����^}!��oi%Z\g���GX�f�~2��?��
:���,�U�k`6���͓�K$�4�+�y���|�1���v=�BM���׎��Rv��'�V�5�v8�^/��뢋��o	Z�E?��8@'X��tj����/�<,g�R�����&6VѼ�PP�XQ���/�x�Ғ/�w��<�(e��k�[Vwt��Q�E���O+�zOD|��{�!\��@҃�;�W{��Χ+�I���LLG�x�c�rr��nl�v��Z!+�1dc����ؐH��f�E?�"�7q��>�.�w}���tAs�)��h1]�e󸱪�n�
�-��0��Y���.)-����s')��vss���K`��p�>��Uq������)t����'Om�������y�ٸ&I���"z0����f������!z&��5�����j��W+2J��l��Ӵ��$�u+>[2.W���WDDA8N�σ�}e<V�w%R4������K��K��L��܆�@�w#Oɾqt�g���Q������%%r��Z�f�S�������S����ڬ!�=��ٳ:���,��D-��ªi�Z"�S���T�^��ǝ�`��w=#�OAoxn^#s�F~~���Ƶ�|��d����yP�ׯ_��V�#���V6��UL�,��u�$#EZƻ7��{�I�CЏj��_Xr$�\���r�2��P�l,:�����$$��7]��,+{�]�4�)Uո���WZ���^�g���e��JHH��������t��$1>!��Z:�_+��u�۞ϐ��jH�	&�{�K�1�=f5����~����aQ���c��U{Ru+u�u���;���+-����V��ak9���G��f�V��Pӻ���埁�}L���?8zffyCv{���/�t�`?m��&#�BN����7+ީ7�ݗ�"�W���2��MeH�m���{��u�'.�zߎ�]Pp�<x�5�����D�.��]a=����ZX���	qpPG
?*(���"A�����
��>�ez�5�E�ֶ��T5%�������C�]u���Ga�����Iw�tY�n�߫�(��N6�w�Ք�L���ؤ��,A��o]Ǉx�\��S%>��U��|(�7 �W�Y'��C�������9��c\I�T#��
ry�x;.T��̓k�T@�f>#��F�S���i!Ӎ6���=R��3d��m�}�܆�	ܳPoMS��Ȍ.�a�	�R�fqe��x�2�k'!�-/�5��M?�����>)웣�M+g���Y>;
J�y��$�KJ��LUk[xo^6}Ğծ�6���w����f�.m9�b���MQ[~��?�Y!ن[��ͪ�������:88t}�ٵ,3�4b4����(F���N扬��½�=��Y����}r���d�Y�(ſb�����0�`�#k}����D��m�-����g?�,����DҴO��Il8��cғ[Kw�m�d@F��5PS�D��Y@a�im�¡�0��݅!0MJ���o��q���W��$��_+{�&��[so�h���[�a�|IS�����n�����Ţ1�Q��@N�՜�;�v��m$0�����n[���Ũ�O�lb������
Ί�`um�ik1{\�d$y�ƺ`�f1tl����C�ѕ�iis�U�p�l������O?��$N0�����w��[ EKs*�Z�O�C����g�����kMG��?��5O�c�DFh��$+�O�,A~�����|Iܖ� 1df6��/��A��Kxy9�ru͞��R�a4Z�ŵ������u���,�J��*oH������͹�K,cO>4�	�\o�������C����$h���@��k���?�hټ�"����\$�}C_�)�d6(�Ӓ��3*��Ug�`��i�P��zmw��QG>�/@�0%L�A
�hd�L�����Ɋ+��R��a�}v� e%cWe�,p�^�"�Ą�i��um1��yL�gܮ���Uz��<?|D}���s
Q��M�͔�D���/�`V[�Y���H!���������������,(�{U��Ƨ=/�Wr	�T/�e2���%��ɧ��^i�OjHP����K�8C>[_h�%�V#����Zl�	1���ے��K��m���y:du�	��'�e7:~���zC���f�e�I#���jl��J�"-�o���wG>��}��J0㔾�⢢���x��
�s�u�<�*���Ж$I��yQ��ڶ@�����6p��\�|@}@����TnZ5y���?��f,a)�/>X�ӝYBdPb���=I�p��n�"�첆�����miּ��xI�TQ�ܼ�$d�.Q&N0�J{��.���F����o�#�����t�~�IAE�8{U;'��#H�
'������p�q'�=��%,��U�>�~�b�07D�'�t���l;��e5_d̹75�$�H�R�I�ڹk��< '?������-���6�8HO��V��>�"�΍�-�~Y �f��><-�ϴ,�]k̢��~���ն����,��A�y���� �l]�O�ڢ�2���5��h�<�$��sf��)'�f�9~gM���X�@͇���q]�*innn���t��T�4��^�^b�N|0c�����ּ���m��2{��$�`�~�?��m�#����@�ϕ�Z0%�PIC�����o�?B��MW ����ϟ?�= ���F��Ma��4��G���=��ĭEЯ�hğ��֮]�[]n�K�[*�bP������0�o�lk۴I�~/݅6��NUb=8�$�؝ʰA�6䒞��){N�6�lJ��x[?1��l�y9�^?�G?�RI�ܐo��ю*�׆6�d���	��}������999�r�3��H�n��-:�eu�뫤7{`��QCa��t~筛��+�p����C���e�%Ȱ����K��FM)��M����B����l�}�Z���-Z�C��F��"|��Ã���H��y?l�\��
Xd�r�I�ōI�����d�S�Iۥ�����zƺ��J��qEܲڨ���E �^���z��nےrm� Q�v7��Qu��ЊGI��agH��u���2�5�j�SJ �@o'X-�J�a=[1��:�Fc>..t3TYOo���KX��`�_GW.AZhwl�@��	D���v{a�)������|a�\AG��r��T��u����e&'����q@'���ߜ8��I<�%��7����>�+��+���,�|�@!=l1�q����H�����>X����v��"�98�a�n�����b��U��	�s�M�]��B�޸�آ�r��-}��j��.wk�?�;8|Y�3v�d�|���ĥL�j��v�J���ai�b���'�~�\��g"������_3���!�:͔� �u�ј;�q������gR�͕�3���VO
����Jp�b2��f_��[II�����u��n�YX���\m�&d`��)z�G��6�h��΃ccC��`�hq=2^w�F�m��{�`��qcF��"b%v���L�㝴r��^�Q�7����H�~�W݌ٶ�����լ�:���2.L�K/3F��I��^nR�醶��ٰ͆�A�pKLrT�����C�q3v?&&��ٗ��4����3~�˴t��c���w7���W�ףߔS:�׫��7���d��'W����>u�	Yt���揩k,~OM�K3-Z��w� ץ���vf�I$H�!�Xt?Ƃ+rr�l�/ܿbY��ᅼ���`T�ՆF���e���V
a֮���Ϋ�wx��
Ve]n��!v��nnn���:%�(�d�}
��#%��d��'M[���F}�;jh��XQD~�	:3���F����#l�ݥ��#&4u�C\�n����N"�N�+��>�X[47����䍲20u��mmo�Y���~��M����b��&=��݂n�[�/���Fk���C�6��~���8C��b�0h'��D�u �GĘ4Mԙ�ڳ}�L�7��E#�� Q(M���Z|�J!��LY�}�׍�Щ��I�V��b""���J���tdf���p֌�^��\���U�u��0?����M�X��`��da��L���'r44n��}B�l_D^�w�j����	߮�^q݌��w������s5��s�c�n�]�
��M�����2���J@Gȑ~g���P���Y��:�ױo�h��Ou��hڀZ��v��6�y~vX��oG[=M�?��=i���#�8�Pߵ��	���-��(�T���JEV�����&�S��P�
EL���;х?Y�Ǧ�t.l��|�<N?2���G������'����>�c�(	�Ș[QQѿIJJ
͟�OC� i�R����![����r�B��yq6�\�:���������x8���NбC���a�Y-���OL�:��F�4��52�J��"��nsPT%��PV}}}��k���9?+����9��:���p���Y��o�ddǑ��D)6���o�:;,��g��N��f��WX.�O�?+3���ۄG��PW����ҟ	��۷o�<JO��� �����~Y�l�ȂR�C�~|xj6�6���4��S+� ڰs�R����B��e����"�mD��|�?Y��<��x{Vz,`�nW���n��lV3&b�U#Cp�|^ �����B3ӓ����@ɾ�P��]s�39��|�����W7w����S�-��Q�$s�Q֖����au׸XnG�thӗ:�ߝ��'��EE{ܯ3��?`?����7�z�!Ą�<մ�����6�AuPW��>�$����\--n�e��G?n�ǂ��.uo�"�1(S��5i~c��������e[��`�!�ww�����%X�݃��5�����]��9�>������R�j����%mL�`����I�SxFJ��%��o�M_�ڹ��� �ʻy)�)�	ߗ�
4����`dFg&e.�����,@|
� �o�Ϧ��衉аhBX�|*�Xe����d��d�����h�wG�>Ii�g��(�$32{�Ӎ�b�Z'ٵ~���'�<xz�z����2*���i9�i�}�X���RX�9��ֻ�y�� ˾��kzIn�?�ok�_�⳵�9��j��o
jG{�����Q�����Q6��qӹJm��!�ڟ~��7qY���K�r����^Ce�]��.~q�,�@l_33�
�%��2rx�ѫ�9|�B�,|�4����v�_j.����
����|p���m�/��g�}��r/r-�Gs�96���T�௺��#��k������?ݥ<�����}��ʚV�F�x��`��Gp���\����mmތ��O{� B���$L�����~ݮX�y���|�r.-���_yfs��v744�w�T�B�����i��Gům%�k�&��˪v�����vԞQ��g�~�N��Ym��/y���H}#>���x�XX4�^��ު�i8ƻ�����SY�XU�h�/S\�����&� ����͚z���ק�������I!~Ʒ� ��~��]D!Y����: )�p|o��`%$8�:,���\<Y��V�!%,�������d	��Y .=��~��Y<#�?ߟ�?�Ll���{1L&������|�L�J��	�4�hȵZ{��(��� ������y��L��o�J�g�e�nY��V���nqRj��6�����.��=�,�ߓ���P��s���=�Ų!��7��zӶ�C1��%�_w]v��@��on����υl`6�%6��0��_K�QL�����_H��A\R>��}~����c+���΀a����>��H�~.�,��JY�}��_2F�1��v��᠗3IZ�c���e��%���\��ۻ�j=�;��j� ϸ��v�9"�ƀ5;;�z04�9�����5$��m��>Δ��z��_J�ytcO��������u�%Wk9I5O��/L[Fd�+o%_X���y����$��{ڋ6έV�(�cii����u;Z��L�r\cҜ� i���taΧ[�aP��@� >CA������&Yn2�
k��<hhp�R~�x��o����l�a�śrWo��_�mn�{���Y�X�Mv���H�Fo�u��p��K[ݤ��=�}8���|��}�O
�,b}�����;wʩb(��s�`�L}$�W+V �2��O���6�5/��YY��z�����˝��I�ď��&���Ȋ���b��?�N�yKig{?+�]���隸b���KA�6O�#5��DvQ�ny�`�mȓa�U'+#c�C�q����S���9G�!�:);At!��YE��</���x�Z�����ٳ������p �yw��GX�"�~!��\|�N���"�.�\��1��|����H���O�կ�9��}}�� ]K^{0a� |w8�����8���R6$�IO��ǅ��Egh���p���mW���'3�U����2�U���%��ۣ? T������,_��������})�I�=x*<fhᬠ�"��'R����+V���b�uS��g�t"eˊ) !/���'>��ܜ;ޟ��l���#��#2c6StM��ި~~��$^�~8��fZ�k�ƛ��
 �}�t���k(�"� 0@�ˉA�W0�P�as~� 5p�+277'U�ߒd�yLS]z���]d8B�]�2c�>l�/d����u$c���_p*e���	�2��M�g� 	��3�Z!�8�t�Y�aʦ(�b����;��p@A�F���.�c&�ňVH�ř6��4`2�B�0�z}�o���\OT^Zh�q�@��.������qV�l}��b���D�+P�����:����<�����+��t��"fԡ�g���hk�aC�	��8�a�������:%\�{�>��=<����|��� ����݄��$���N�&yu
�i�+5��)���G�)P��lȂ��m��D�*LT��Ëf�=6`��-0Z�r�*˯<��R�N�C����{MD�>������G��Bډ�{�H�x�<6V���ͶJ�������Lf�:·��s$sii�a�c_L�IH�R����B�7�=�$n>�"�b�$xRq2wJQ哣�ε��&@J��z��ӫ5UW!/��ydW�Dwp��Q�x�!��9w*��׀@�8^���ڎ>�t ��Rm#�`��ϱ��?���M٪?��عn`�{P.�{w3y)��p�bT�]��^���)�WV���BֽC�^��B�'��r��3��as6>*�"��b�"u�.�s������鷟R�i��0r^|o_�vbeG�%;�ح�E����ԏ() �'&��1���(F-��@��.�u�O=v�vv��<4�������_t,��r�v��^&� �y��~�*y��u��I��<6�r}2�I�	H�n��p�B�� i _o�B�?��,����m�I��M�3��&�!-��� xh�䉽�>�3wyY�O.,�B�޲�n��f�%|~~��	����O�.q�@~V4d|� ^"���~�@�4���ibe�4}����
	S�ɥ�.'h���gp�b.胣06��7�_���j}���k����|����o�um��H�V��*����$1o��E���BΛ'b�|H��X�ss�8\��Ww�Z�i�$��'�8)P��F�V9�\[�B �[�ȳ�s�������s�Yb=_�!���( �AZ�6�[6"ñu����4ֆ�Ho0�i�@���4�5:�n�&���,Q��'}�[�!A��U�x�J� w�W�{�pъh��N�S��xYL��p������1+B��**mɰ��'��7�l��Z��S�tLo��Qٱ�۽;T��22&�!���W[r}��Y��G��S�,��(�|��B𙋆Qp�+��@.������C�:��6S),8g)�Vk�ģ�5Y,���8���W���A۱�S_:h��:��|bI�S�D!LcS��pة���O"�?�L��H5Q:xx���j�l|�'	���چp��Y��J�� �#��^ؤ���gDV撣��UG�	gLYV� n(��_�L�M�YN��9� ��U����<�;O�|�"�)�1��"�r�h�ρ��j���iE�тm$���1�[S���0�52��nܚ&�,^�Ű���]Ŏ+�Y�Z�8�}R�.�%ӎ����*�Ǣ��G���`<�r�{���� ��ڣ�K�j�Y�8T�gC��9��i������_I(����d�|7Ok�4�� 8d�u���͆*t��
8����R[�E������xz�DO�^�w7�*�bއ	e�����jPb"�L�\��NE��{�o�j-��@EW�t���7����x��E0F�<��Ä80v ��?��r�ڏI�Ӟng�6rZ�E�^�¿��r���0è�F�&��՚��`�a��kI�Y�o���4�*_��H�Y)�o��2�w�<����ϸ^Tϔ5�b:�{� �._zX�V�L�����S�o$��톱�bIa�Rڬ��3��YIA�
�.*.�eWԲcR�É]iH��b�v0�v�~����`����*@�=�XӼ@�ᐴɹ�,����d2��FM�SBV�4��6LaV�!a(�n٩�k�w��$��8��},���XW�����uD!5�)�2e�fjɴ�O�h��(���o���<۩ѸV�-���������
j�Ӳ��'�?}���DH�g��6��d�9�f۹�$e���%���j/��X�#)��jbc��Y�|�K]��p�
TG�6L��Oax�I�q�����3#�ON�^��ޙ��}��3r������;���F����z�Z��,6]��K/���U�,14o��Pra��3E��>�H7;?�ry����n�N�a;Ѷu0M��2��h%`��1�
��r=��u�߫��.�����w����]�;�0�Ϸ�3MO��LP	�;L%yeW:���ܳnѤWRe�-f1���jۧ���h'��&M߇/�9����y,�K�Ll�=��1Q@㧶Z	�{��D|@9o����[�����)@�͕��4����4���r5v,��ϰ؏{��,��Y�����J�3)-�[f{=,���,�(o6�i#k�b��Q��V2B�������	�َ��'X1$��r�`_�cI���â�E9hU���,��u��q^~-�'¯y�GH���'>����Vdx<s%UH{�(���#y|����1X���	^����&ӝr:Q�r�D( H����O/齆���B����[BԉV�А��:/�C7_t@o����Ch�t��o�A+hnG-�?i��{���G=.�ċz
wٹ��t?}ș�=+���@��߱��î�H*'m�12��ܧM�ƗI����+�� F6�¬�xb9��~zjz�Ư9t�^����3r�����bb�q�a�a*N8��V;�����ō����F�*�h�eۯfp����X��PA�';�&���u�6B8���lM����lܝ:s�:�6z�A���=�gm���v�G�:����=rC�%�i���4޼3��+�9C}ƪ����7�S�Į��!D�~Oq`g>፞ܧ`�j҈�ND�gL�D�T��O�Z�$�*�E��k��Ğ�2��y��=q��y�#�
l<���0������)qw�߫Ʉɴ=�o�Ӏ2+鯱��Kz��8�ݛk��^2���܋��P�D^=�;�S~�l����o`
�lkbB~x/��W�d$^*y�X�q��V���!���Az�}{n�Ǟ��-���"f�ɲZ;�1�
��d��T������c��1jd�IHټ}�Q�P⟠ڈ'f�],j������朋�(�p����I���Q~l���Q�7�G�Y|��}�k�����_�K�?Ў�B�1���'�x�閖^wT�e�����|�seN���WB&{P���QSX|wȝ�{F��ٳ���n��J3��]3��_�l���y��h���SUv'���l���2��^Y��Ǎc�oQ�O- ��HgQ�P�
�Y-P�h��Ui?�S�T�~��P��U������*���NG����яm0믣t���:8T�j�(��0�T��,��\�,�����=�rm�)ɠ hɲ>B�+WfQ� b�z�>���b���%h�F����A�;�N�e�lh��!~��̗*2�����sC��6�]�'#�z�N��҆>F*Ά��N ��������[1�q����QQw�y�&��@��g\�*��P{��o,��bC�v˧�5T^�a`��Z�:s�l���q��Ն��J+Ͱ��OL�0��W)1Qs��Olj���>����0i�X�F~f*u[�-:�
�4Xp��4"k�,%�Ԋ�<ğ�G�h�"���H���e�b��+�!�ߊm�,�r��$З<9zU��N�<����N��p���VJ�:n��(:(U����K1�^��R�!�r�M��$�:|�o(�?�WޖP�鷗Q�t����n+�6��=�k�C�3��1�+W�I��R���)�)���V�G�7��.he�:{��~S\������*|�I	�Y��!��(?�/���S<X�͚��10��9#�>��ۯ-��� xG6��&Sssu]MJ����{�ܤ�'�`��Iv� �B^����'xҨo/3�B&���c����6���r�5J^и1�=��3<�Z?����]�P"�.��N��K��Z=����ݾ��5>:*%R��S,?b�>���p�a9�<�O
ކ� Ȝi�I�촢9�4��&��h������tA7�F��|��ܑ9_rY0��dsY��j�0���J�Q�"Pt4�</U��S����nu��R�����_�͵�)!2�R��L+���}sp˪u�������W�s� �`�f��UrĿ���C��Hџ��Nm�O���&@��j�ז1)>	NT{��܀]�4�� �P������#���⃞u��`�%?�UV�+��r�4e�wN�w����+��Q A[�K�t�s�e�Qı]]'n�B��eH�WLz?�����;�Ֆ@iG���)��h�L絃���ec3b�]�
�bG
���~j%��s��s�t���bL�d���z	�Dy�Vf��;�T
��3�ݡ�Q�-S�'Q��?���44���,�x�k��3W�~� ,ҢG�ĥE	����YH�*>�&����PЯٞ�͙H�'���F@��@�O��Z�3׫'G�����8��[�+��T/�KL�����h��)퍖V����-D�L���4�'��s{��]8���!$����;���B�� ����?�����U☱�+�&���䷻���[&�r���/��`r[ɬ����Q\؏��F?�ytW�b#.��[<�@h��3Z3>�<D��p�rХ�{G��������0�Fi�3bA�t>��n�(]�(s�&�Tc��7�²�������s��G��i���e�L1�����-�����x7�3�Ї��w���Z�� �u+�ڕ0�7�d&8����Bd�����|��a�[q�&�p��jFR������>��m��E�X��ZĘ�Z+϶2�`�B.U�<m���ï$��m���U�
3����,�+=�H�-�	YJ�5����ZA|���c2�Ad�aB��ֈ�	�L3�	�U(�B�LI�M|<�	U��O����sݬ	����	�90���Z9_�8�9�S�VpMM;J1��3v���]�>"��?��Wy��em6~I�� ���(f�&��z�
�]������$��y�,��0����P����d�ߤ���L�I?d���DF��c��/?����X��TڜMp��ͬ����h5y�D�Zs�́�f��$OG�#��H�b�t'�Q���5��i��<�UAs$���*}}��.�)���tđd����Qj�`��yZ��Vf]��5r�R�QLr�ՎJTfӷ{��>��ֺ�r��U!ɔ�"NE��Q���&EI�~���p��lѪ=G"�eumJ'X?�#K��٬���:R��>�oB%���'�AZ���v+N���VܻnNI�.0��E��Y��q���+#�������u٥�y;�Ư�-?~כ��ݪ��ڪ�Ym���i"pyV����Ƚ]<%?r�}�Ht;��|��-i�cޠ?��΃j�̭�ӫAv��f]��H��;���G���GQR�&�u� ʿ��j�cJQ�p���l�G���л����l�m&/��9"�ۙ�P笶"h�f\�j/�<2����.{��H"P��V���e���E���&}�L�F^���BE�BrN����W���*[�0�ù��B�O��rr��m��P���d*��?e�C����V����x�z������s8z"��O�vڰr���̔>2��?�V!u��KQʚ�K}�����1/��EGk��h�� �����+
,�~FIP�Z��\\=]L�����nw<�řNѫ��h�2��Oaq��> C>g���r��w�l5v?k�-8\Cj���LՖ��s3$~�n�y�p�]R�3liL�}��X����Ȣ�ms�KK9N��H���];Z%t$7ˤI+��%^ㄱ37׶��q �vZF�\ٟC�zg�gp�
A&���W�԰����]���d/�5��ǿ� #��e�����P�����9=<��խ�`$�R/L��@�A(�ML�4�䌙�MM�{��j%V[��C��A�A-�p��.�Ο�f�d��q��i�[���@���P��_$�4���\NU6l�)���+B��j9G|^B��&[=h�:.�z�|�M�o��qiҠH�AB]V��/p���G��L�&�F(9����c���8v�i�o+�G�ˠ����cp{���2��]9�g��{�[M�oE�s���Jꡞ��S�nR���$�9j��Y�Ѽ;�L��<'@J��)d
�3�_5��W
Fh��h���0��[��B�Ϧ̯#�O��W���s`��h����������(偻��+��	<:��c�X �z��W��I��h9j�X�)1�u:[F���k8�eq^���9�4Yj�z�E��_�+SBx���b�%�D����Mr}�N��z�{`zj��PXɖ�$)�m<{�JP�`�6 1Q���3 p���:E��������_ B��-������j�W��8�xrB���\k�

���Ey���������K�ќ%��P��da�GR���6��P��u?�*��n�	U��]�6_F�����;��t>/ұ�(`�ذ��ăU���q�̮�T�w�Sqv��f�}��r֦�&"�(�i�	.+!)�����B$���?��6�P�Ô�%-
��:��>�g~�mp�B�:,(%��cQ\2�c�왼O���Y�S�w�Os�d�SXߨ����)m�Mo���煉s�\���00M�z������S����;��J=��E�6��pV�ɈW��U��f��C�%���?e��>�ܞ�Pc�̟�я�����|��E��0�����|�����:�
�k�d��'C��'~3��䜹j-�a���H��O}t��6"%^c%�¾�����a���A���I�ZZ�p!�J���?Qn�j'U��9r��FЂc�:�5�?OJEl�H�f����e&�E�����${�	x,����BP�a�v����	T�p��4M�6G�UXK�>I�Z������K)]aC������kuΈ��ՓC�Ki�WmZ�E(6��G���6ȉ-Y����qn�+����4��9�H�Z$����7;�������Z�F#C������s�Z;{ ��J�)�Ge�g�՗�F��P�k��pqUm���S�͕��[���R#�Q44�M���*��Q�X�'�(!�Fz�+T?@\�zP$e8a� �-i���,%�'%3��>�^�"pC �-�T%㻺�v,��	��*��b��d�Jܮ�{��Q:g+�"�CZ������>��O#�a�Z��z^4�����#�G��r����]
�G8f�lt���jx��Ѩ�yC:nx�f�/�}�����������կdµ/]����ް;3��Z!j�*�A+��S��ן�<P����#
\�]S9L���X��<������|d�����]����i��h��߿�O����vV����d{7�j^g����E�H�ӄ�����m��ᬥ�_�z�ו̣x�~��?G�A$�ځ�L'z4�~/Z3�D���Plb4Cqn >���ݙ��?�������n�V~\�xx����$�4�P�b�����zu4����^o� �$^b�~�^��Ň�#��;��C@(�b!2;��\�g���m�d�@���oֱ��:��0)�R^���%�-n>���v��x9�P�y��Z;� 	�g�Ե���F��>)?���y�c̼ǆ��\.�Q�{qY(L�$|�����/2�7�ebP~�Y��ٻ�0���*�.�q|�+�!U�a��Ʋ�4T��}oE%�aջU�Heև������t��#	�Q����s
}:�NY����[�lS,1,gT��)e+u��-����K�tb�Z-�3Mj�k���ҵ�P������$���n�G�� Հ+��d�����/�">1�S�BK���a�Ň��X�F��;�~<�JӀ���c��45�xy40�=����G��{�d>�A� <���V�Nv�)��re��i�ϟ����¯����f�H:��P ��B�ʗ�����ÏU��4s�dTJʊ�r��������"< �Q�KU�d�ƹ��kg������Y��g��~uM��(�*Js5�h6Ɂ���X���'���֍�(��������s}_�!KŰ��Hd���rM�'�����F?T�vr�h5��{� 	�^_Y4t�1 �)r�����x��]�*q��}���)|o� ]Ʒ���Ix��Ô�̷�������,��)���hv��`�c1<����j���}�4���cF{_�#$zat$-Gm��f����6R�neJD����.s1m�'��U)At �	�g'��$ w�B���?�������=�q$�~��u�>���X��׉�aq��մy)������]�9-�V�=�s���X�X�T�Tp �a$#bJ�!܅,�T��FM�W�򭾫�@κ;R���R��\jq�k����	��V,������W(�I���Iw7�飃QV���u1�����۰m���E��9�1�����Re��#����@8�A�H�s=���h}��e�[hh�լe�1}0|���Xe�?�ՕоÞ�l>9����
^�BߠyZ��q<���83�3���]�����7��!]�V%F�1���vz��_}:�<�ލr�1z����"���xhV�g4��:��&��M���t�@(>7l�~z{	hVv�/����8��/��+��J��8U	�KO���M�%�=�~w����h��cjN%��i�|���sݱ#�$�98 ���� �tzp�Nm+�0QU���e�Vle��¿��>�V"��Aaa��!x���VhŁ���قLB�UFJj�U	���Y9�L�N�D�,ӷka���7�)�^/-߷o��r�klMObUY���A�4�Ph���>f���n�u㚰=8�"�?8�:���S�S��>��=�iF�G9U��]5��%�W��#�ǒ!�e�勺�(���CpḤ�á^6�Q��Ҷ���x���������J�W�4��U�Ϗ�Lv.6k �sp׀���D��V���I�Knw�^Ύ�Q�#&�V�_���$������mH��ݳ�f�3�~Ek��&�D�q����=����+������ż�4�(}h���Ry4��92��_f�-��J����s����/���G�{����ZVH@��ɍ3Sܹy��J�e������zSd�� L��f��X(�p�1c� q]��]��BTJĊ���\Cp�e���0�0 @��;:*��O3�P�]��Id�s������|����$��\�V�ň���[���'��|%� ���<~������z�I������؀(�_�M����/g�YE��w|<%b�����uD��Zv�D��Vo�6|s�$IVU���y&�pw��V��JH����������j�Uy���-R^���rnn�V)�3�z��տ�[��η���<;���7��8���w0�p�Օ�兽Z��ɨ��F�ֆH	�3��o�o>(����'�[E�T�H��e�2�b����o&66�>C��c8��"�u!���_��{�>g����#49����;���{���k�+^��7wR�2����}M�/|e8��f0��X��7��_!Fz7�Gޮ2���ԥ56������&LdW�� 4[Z�����UXֲ�g���p�@��g��ͼP"49С���;jc�6�iOp\r���c��Y}"�r������*!�!t�XM�ȇ�ˡ���N)`�Q�B3�aAl��ߍ���6��b�.���@�2j��tح�mKq���\]Z5ƿ~X8�TTdS�Ru�)�M��A@�F$���Um}\�T���i^�2W�� <�fϩ����;Q�, ���V��AutdNKKKr��A��Az���|��g��C�uv�� ��EH�ӓ��"Ne�ds��2����~��I�~���q֞��@��1zP�8/�W�U�O�>h����G���	V�KA���j������ࢢ��v&�2u��o�H������\�2S��Pl�߳���H ��9dM��H��C���&���/�����4�dbf�a��ߠ/���E��41�- rB �m�?�q۳܏��X���2���C��q�}��¼�+�X.������{t��Mϋo�A99B~�\�C��3%�D<,x��c��]O�B9��U�L'WMM\M��J��p��ٓ��ѣd�H��#�M��>�f��ɿ	B�|>��
���{_o���^ڐqY���3`[��}�J&'����0��Ź��2c�8�eK�����EI�N
�nZ
�qD�^�z{�F�2����(���SQQ�-7ك��u�[�,�q&��B�I�-fʶi�2���M.�����܋]~��X��D����U>�v�������o�wz�Н5S} f��~+�*�ܜ��ϳ@6��m��'��#^��_��$(��@�9�!�����4��*�O>���J�
�4w�"!Iη����d�s������.t�ч��px���m�52W�y݋l���{pk���ɼ�p*:::*#''V�>������u�Iv�9O��������յ���ǦQI�@OOAJ��݉��z��RIUS���41�۫���^e�f� ���9q!s�'�Æ_�R�q-�sΒ�����3�����8��3A�~�r�Qɑj2a���YȜi�u�-��w��dV�X+ؿ�f��MGˬ���@�h ��\�:�ڎ�Q�-��i��e�g8��5���W^�)IZ����1?J��m�+'��X?�:Ŀ��ΠxJ�ɒ�5� ���?d7Ԣ3�ׄv�5��tک��N�d�"�u���?(��� ��� ���"f�Oj|V�Y��f�7eC��4lq==���ְ�]�j��,"vk����ŽB�?�T��\��#:�1t��p�HQ���nu!G���?���4�ĩ�/��d6L��0�~b��n4���mR�+�˭�N9���\��6�x�++�g���������Sz:FƬI 
ژ�#���'�'�O��ogW�?�5�Q"� G�_��/gԔ7Q�5&�/ʔ���z�dML�=W�q�=N>���/��SH{=����o �l��C}}}��~a𶰒��n���ㄧ����y��ގ쵲�&t쪎�N`|vF��X�u�z��g�5p�!X`,��j�S�Kbm��e��S�%�����r�K�I��$D�e}��}�VT�����a8;����oo	��F-�v[(�΀!�]w}���@�aJ����4��%��}�}�C*�Hh�#��t3�ʟ*�[���@üۼ{��v7� �M:Z��1�M�x
 xo�(J���O��s���X�_r�ಝ.p�U�P��yv-
`_l�����6W��ghB�<{�t�r^�g���a��~G�,$�)���`ߣthl|GR��H˵ʺO?�����#�{i�?�O+��-������G�g�	��n����(�1Mx� ��pߗ�h���%��f�/��=�4N�a�����{�\� �	<�\T-;��6��>J�.�JL�����i�-D��h�+��[t�̰�e��݋�����M�u��.�Q`u���z���E����� ^�`�2'��y\}uc.Y����c6vɶg=���IN2���~�������������>#��7���*����o'�K0�����ǣ��r��T���Px(ﷶ���Wݰb��Z&!��|��}�@��_����A�b2C��BvN�5����RI�_�����e���Y��Sfw0(�����h@�=�o�]#�����H�VT:�\L�WA��PM��#�SX���3��o�O��7�'�}Ū��#	=a�!iY"D�*��������g�\m�X���x�2�O�����J2`S��[S܃M�u����3���(k�񿧜��䏹��bRg�j	�e
]#���KF[�$��(�:��a:�7��N�RJ|��l1Vd���Ƒ�Bj�O+&���0um	��:����N#���X��O��Xq�	���]�N6)��_��p�ܻK�2��&����#.D�4N{��"�,�Gd&�},�q*�Bnghc-���n�I��7�y�
��������~�����l�%=�����d:�wC�?�K%U�q�\�d��)�E�͝ZXXv|s3�B�j6gw5%��i��U�ꑾUA��V��oV�dˬ�!qD��{��<�(�1�!43P}�"[��:��{|�>0�;}9%�~�O�v�
��z��/B�A?��=j]��6טZv�������,��2�A!A��W�̾?�^�ngԶ�g�� �wb����Bϟ�A��o�g���B	<�$ڭ�%Wwgon�
�tJ��;0��������ԇ�7Bp a�[��á�P�㽥u����N
����dҼ����y�lu�Y�!��)�!�׹֋���Պ�Pw��A��.�?E+�]aXi�}�w5�V��D��
����p�r���L ���Is^.�?l�^�"�{�P=<dǌ�=��5�N�z+B��]y��?j���˶*������UǑ܏GUr��K)�M�p���_��\�Ys��C4��A5z�m/ŝ��aK�����D�����AL��f΄2�hy,�����k��F�jc�[Id�?/έ>��s���U=��o�J?ac%���FZJi�8�l%݅�LҬ�="ݘ�rsRB��[�a�l�a��-+o+$�� ^��U�Ad2<��Hi2�Z�������𪭪����[�o7���%����Z�Z�Z�kX!f��l},�@HB_7`�ό��q��0Ѭn���rm�Oi�cQb}Bw���2G������!6��xS2�8[��c�aE�8883��4\h���н:��o�9B���W:��>�G�3<N��� q	�-��1w�[�L	
khh44�n��,*����y�ԣ;�e���&����q�����~��
L&�Q `(���x(�1W�v��e�����bU���Zfl��)�7��	?�(�+� 1��%F�^���&��:�Mݵ���	�Ǳ�Y<�>nx�y5Z��w����5�>�|��Vc���(�H����_�єfƵ�C$~1��:N�x+V&*y�|VE�W5M�mw��txť
�+q,f9��WN�wo�z�:��s��A��~Z���xm��H�[��pA����
lPGi>�J��Lm�;j� @�+Z`2lS���c��C�釼�ҮH���kttCy�C$C������p"~���O��^x��? ����8�t���iR�H5'O�m�GS[=y�hob�����b�uj��@�D��zh��O1ʵ����{{g�W9&�9���"`�4�.�Wݱ��͇S$�V��o��7e��~��Y��bu w`�u���|���1l�����#D�x����������aUn��Z�o=�yuVI��EX�_��?��00|N�"�У6e�����h����5��5o�y�EY�3���"��+��h�������AN�J���L��jj}S_ܤXq奥��=��N�h�6_I_��T����R���./7�(QӖ������F�ۭ5ԉ���I/݊��}�{ު�=���s.�_�SR>����h�,�(�<� 3�S%��;Y�կ��bH'H���X�����4Ҩ�����$�f�����z5�;3.s���� ��;y�3S羿r|}f�=�Q)���*eԾB2��S�7�J�ӝ�D���s��Iq�j�KD돀��И�i��ah}�F7T�M<�V�MI�J��I���d��$��x�~v�Y�uS����յc��W������Aj+�v�È���鉪2��{��.��3�/�q��9X9����]�Ā�ʱm�A����u������C�����It��_�)]�ry�Io@��S2���t^5�%�>�W�P�B݁S���ǝ��;�T8IS8�ť�m=��"��A��� �h� �{%����-��p�����{{k�
�����h�~��!�S	�0u� ,of�娮ZZ�_����(��=
��\}B�,S���-���[l�S	x���_�g%����M��TVF��m&�mll�[�ʚ�Q��23�YD��Q-�i��.(*
�y��6����]� ���_��v+-��w�v�{��[���ui7#C7��ԇ�33��m��zqDA���Ge��?� �bȄ̙�@E�??R3�C!aA+�����Q���e�D__�[}=4�^o�Q�p�ש��4Q��0���WR��/{�LH�:�Of~�5�D&��_�Ц���Sg4����I�ǩ�>�qi���ԧK�c���3}�!���2�����:4U�{��0�$K����.Q��>^���P��W�ʓQL��~1�	_B� Ar��@��~�l5��Q�C�s��d��`@��>8���湉�BpZƲ;Y��B�w�}j�qS��(���j�O?#�#Q�.F��������vF���N����9��v8T�%���>���IL
8�G������^������&<��|?����w�+q��/x;��PP�����n/�u߉�P|�kna��M�;^�ݝ����;bP�����q��h{l�S!���ħco�v������ݩq���l��r]7��U1��K��LHf�
�}��I���]���J4o� �؉��&�Mk+R$��f�t�FU%�?����u�ޞ2L�L��σ����}\4C��5�+=�ˍ���L&Wྫb#�F��0�3c6LE�m��C6�]�,����_7��Em�0� � IpA<�'��%0ww��\�A���[��w�]�����{�U�GS�{V�e׵��^o�Mq����$X�{�~aD,�V`�β�yv����ZX��w�(.7uS*�x���?$zMz�Pn��]�qp��H��=�-YBP���5#�Ͷ��E��>����"�G��;�A�����O�xH�JW
Ͽ#q��t���Kd�ڸ<�ăG����w�[��؊g�``aD˅=@��#�a�[�)�yvB�><�1>�S��F�]H��gx��؟]��x5?������"q�FRSW�Ҹ��x�{�5��"���O��uS�$9�ڐ.�S(]H㳷c�����P�׭=7� ��r������u5���$�,,���`
���B3�ï$�K.�3Q^���ޯol�|�ǉ������������������[��Z���FY�Q�f9��3�u=I�ѕ��[f�	yz����iXDR#Z v��7�M�&N�������(C�F�-�&w����YJ�;��*P;j��&xh-*��5�p���;?�o�=�HR��&����$oLC��|���)a��7tTj,��'gM���v6e��ETF7-^�i����TvX�2��︔[�g E�x�?f/AO ]^�����Pޢ� ��l�+�,�1�!M�k�)ng���m���Rf����sU�;tC��h�h0���,IW2ع�͠��mڊݧ�	='���J�+
�e:�W��n��
�c�����r�H�P<��[�xF56477W�=?E`��-J�n?�[��L3f���E����bH�{kkK�a�����78(����HS/Ta���%K���v�J�D�|;l�p�,��,�Q�zd��,�Y4PX�@���\
��mh�`7�dL�!N�����I��#e���DF���TR���{ P�y�Vk��טOG��N�`\e�����]@�o����p���v���`;�>G���xE9+I�[�����W��2YhpY�
�G�蓅6Ѥ#C��T�숾8�k���� ��1�e��[V�*^�wm2V�C�4/,[:��5��IJ�!Ɉ��b���G��όmw2�+X3^e�K�� ���7���Ɔ�z	Qi�<^V�l�=ܞ��9�'1��L*�x�֕��zP�͏���~�U���n���#���R�nY3��it���Q�0����i?��,[�<~��%K����K�ۚ����e����88��������ZX0�U��$�+&%EZZ�<:�疀���A�ۇ3S��߿���D�&g§--p����U:�+g,�i�!���#��5�~��"KA���95�*�lR���A	�T2�&Y���;p~���\2�ch��=��km��ݛ�oF�RUpH���w�H5�ZX�`|��zh�)b��Sv�Z;|x"Xé=�{�:��Al��~��<ϡ����8L:w씔o��)����ϵk����7I�W��N
!�^e���VK�e �v�I�C�>����Hᄑ�g�<$�J�p9�&1A.M�/Ҭ�Aȍ��ٟ.4ߴ�O�G}�UyMз��OO�|�%//O��ϯ�|��Einn����Ҽ��$:<W�����B����iN�����,���3Eޫ��D	|�fɸ�54^�����Wӽ���8����|�;����sp�����t�F��e<�H> �N�/>m��ᇤ�g%'Vu�'�*�n�)sN>P4�QÉw�o���}�43S�����r�-����Ʀ&`/g���S_�1z���n�v���➔�x1ܜw a�T���	��q%��3Sھ� `xR��s��AEy��X�ZYy�5�nnE>[9�Rd	E�
�+s	��P�/������q�iSa�p�X�Y/�4���fJ��4(2�L�V�m���gy~��`>�k��A6��q�	�u�U�g;w���r�>w0X����������j�<1\GM�5Uz�E���-b⹭1�%�0��EN?y���,ޤK���&Qچl�]�`�NmW���������b7�g9A�p�V �	�ӿ7]|�N�D�{��=%����������Ov��]�g��#~��3����!�K�b�^U�8mzy�Wh4~�K4Բ"�,��4�E^XVT�4KD{'8ii���o)1�dy_*u��h��Ye���L��խv˂����D�KR�?������=vw��ti���%p�����i��p�F>�q�)"}u֝��J]W����9��fs�� �����\��A����`���j�/o�4YЃ�����w���Y�p��hD���ׅ�L�.���m>_���>#�i\"��~�_dZ��|8/ni���y���w9ڼ��)����1=����1//�V� �#ꡁ����>���م��
��ѿ��r��� z�I(jp���b=;����i��Ԋ�Z4�X�e]�����iM�ȯy�z`O�5;���4��Ϯ�����G�#�C����螇ul\fÄ́ߦ|�1}S��>UG�^���	K��2H��.�[���f,ژa�:��w֘�>�!�������M���|01���d�ҡ{�>���")¯��a�h3�R낛d儳�Qe�&���%f�u=R3���}�~���g�̾o@���T��r�2>)ir�x^�F\�br���O�g<za7g�<S���G�a�P'�YB�*z�"�*���۹[y΅�&��5bL�$�u=q>.�ϨD���%�w�r�wYnq���x�ʮ��,jm�LD��\W_�lll�A�.N�:�G�����m���FA�����U^��/���_��Z�5Jhɂ��+��g�oF�������G���|���A�����|�v�:�_���/�{J��$-}(H��G*\��{ˮ< ��b�XI�QR�3���#h sCC�N���ݴ9�|����τp���;BS��J�2.�� ��*WI�j�qs\�"�d�w�� �F`~d-�t���i>���vc�Aϝ0,�\�Z�z<w�3�ܜ4<H��Ǻ~��cN,���"`0�������S�25����c�9|=�S g�``�]���N̻{�kD�87&n���պd�=+�-`?�ȉ������>jo�N�$Z�Jpkq���w=��6����%V�m%%Q���qq#l(�TU�����Q5�W_��Qv��1G�w�J?ش��	?�%��K6Z�ju>nm�F�.��<�.�X��@E"Gow"�r��)e�ٙ=s��W��-��
ԟ��C�v��8���0����oD��X`K,������>�CZ��?7	8���Mb�ҩ���H�����K�}��;?m�J$���J�Å1����#���(.�ORߙ��C�?�x-ݍ�e�ǟI+̘�T���FT`Uy�ɰP�����Ȣv��v̜#G���>���&ݵ�S�W��!-���K���� Ӄ0����-!�L��x�֤�Uq�wj�w�	�|�2��y��_�ΙQAW���L3�,]����\$Π���d���wW�:s�5:���!�n��ץ;���-i�O��賻���$q��
(�vw�����s����O��q#��Ty2/2�ݒ�����%b���	E�Kߊ�'�P4�j���ʾ,}�F���>�cgǩ�QO�+�i6��x���c����`O -�EG'�|ϥ/s<�T�#��\�N�xNn��5�~ge"���`TV��HN`��Y���dLn�/붨��HG����%R����=ܜ�.��#2k9���7\ly>�a'r�R-�;1�R��	��ڗCI��hpiɟo��g�Y7��2/io��k,�fn/���0���ϲm�[/�S�����U�ZK�0{/�gƴ���X
Z���<��Ƽh���|w��	�jqG��V�Y��L��|����=v�0=G[F�Y��;8<��^��o�sŔ�}���sWv�Z�k������kLss+��~� ��	.�XQ�e����>�� �MY��5���3�F	�3��	��a`�]/!���E~�?�)fS��˳��D))�,���z����TKqi��,4uR!�b�����X�EƘ[`thhVCC�����s�g���/�����ud�&v�00Q|�.��c���L��|��O ���+w�7�\�o�hd?d�OLVj��6���<�BE557=�5*|�y6�M!pv��E-5�O�RR�ML(�����9�as�+m^�޷[���s���3p�ܰ�
���u G$dw�V6ѓ��5#-"Bʆ�i���9�dY�����+S�w�=ˑ��d��}����͡a�z>���K�iZ=��$�KT�.֦�<?rJ�0D��wYf���=6Ѝ�Y)���/ȩq���)>�z:��`����/z�^���՝C����"��0�Dd�˧ǂ<Ћr+�#���`,!CI�m҉�H+0�BZ�O�B�w�>~䊀C��41�����8�K�8?S��yڜ��Bj�XdO�?$`c��^u�I"1k�B�����Z�O���/��=ZR�wqG��=!u�s~ibI�L���O�# ��1�>�u��R���?jN���j��?��i�~74���r�e��111M�_.�"5�'��AA�]�_�I�Lou���{z�t@��Y7��/Lsf	���y�ɋ�eT���%���������j^�K@Pm<�Z�T
{k���ى�����ϟ�be�����_zv�R�Y.��zD�!�L�u��Z��cۥ׳"S:���F�My"��cF�Ǿ@�����aG�!:������~b}���Y�NJ�-8ݰ�C!�֩��C�X+���5eO�u�m���u�wqP2SI�������"����ȿtZ�;��W����+=�5��I����]�&8jXl�{���>,��V��ۮ�ӽB+��$.uU�H���,)���I.�a�~Aϐ��a�̶��h`V?_hVug���UT4Us�cR���϶	$�j���C����ڟ���Rĕ9�lx��z8�7�$n���4�hD�"^Z	�4OR4�E�?A��lOc2KM��Dj�t��ŀ��q'&&�`�W���?T���,é���W+��F~۵W�fodh#�A|�F��Gb` PVa<����y�)�C�4�K{^�?��uLJ98�̒9<,goo_ ǆ�koG��isss{z"��%��M<�ڟ#��ީ���$��7G߹TRTyc����j%��Ґ��X��qOaѵ{���(.����H�5�G=K$����b�M9R�?�Id���,���r�5�	k�j�.F������$fR���Q��{�-�g��%�M�[5o9O�_��b��t9/�7B�?�+��=V��E��_}����N��[׏��1*���xǀ�(�s�.|#���~�vg���f�Pus]��oy_E�H�;������($��8&�9�R葾d���&�
��rr¿�Fv׭��t�X��e���u���Bgv�E���+��N�!mx��q�Z�؍�=�{���%��7��VF��"��I?0JX�Vų�s�m`�\̂�?�Rk���
��'Y����������<ϥ����Uo9;�l����0���1�t$[��*�Ƒ�S3֒�Y�o!a�b��Ec�C]ē��R6�PnR�m��q�Ђ�k����M&<�4��Id�����}��&��� �  �X_\ʮ��SH��������w�fk�\�C-X�e�]!NPT����F�t�I3FІ���$@V}�H?�Ax�'V3��'UCȦ�bnD��P��+�>��=ꅨ��~��]?�]-i���ŉUе�u�v���j٩&��~���i��r���+�/��;4��Tn�c+�߷9��<�P��bh�e�h��sˡL�/���<å|��^�O��}k�La����x኏g����8k���nw���[<��%%o�P��,	5�+0��xl����x
<���5��Cx���75��!)�������'�µ�On�a�cc�jDUEEw��?�)<�BCC7ȣ��V���~�u�-6!樬�E��l%�oi�:��ZB�&��O�"���%x��7�}���|��:�� D��}K��ivtJ��ɂc�������t���9@�8��%,�	]���ɢcE9@��{sF<���8�4Tj�yZ����WKƣ���k�_���j�<��w,"�ʝZtP+�Z��@����L}M����gH��^	�
p\J�
Y���7Rt<��� S��#��P�����iR����g��R�9Ec˓8w&C+��� �����9F���p��zjX�[>Ƒ����c��~�^m4�������ps4��6Cc3���{0��uk���gd��;3�НP��=�Y7)+[Sq��h��Y�������`8eW�q��o~�Yۚ���|���I�q����/<gXl�1����B	P��_��2&&J� 9ψqp���8�8;w��4(��Jn�k<�fʔ#>!���|��l����]"1�D��3?��k�H�i\ċi6`¨N�G?��"e�$���j�^/o�>�X�����{:V�B����lB�pq�D0Z�������𐣡}��`o80�o����{ľ�A�ъ X`�"l~���ʸ��Je�48J�6�'�����]hUO�r��9ͫ�u��"c���[��l;�7�_��L�(���>�ڊ���߁=^$ȯ�y��H1�"�<{��qd  �?��ɷ(���Vʽ�a���uTf���A��o�KLM���Q5G����&0W6�AcƵ�tL;�ZYY��%4���\�G݈F����_?�Ӎ��P��-��w��=��%�I�����	��OS2�8�|��칗%{���|�ȡ�����&$���]�ϟ�

����e�S^>�>*���\�8ȣ,�9���x4]�h�>����)�>�=�#�22a�S�P�V��ޮ�|p_�1���R����U������vr���µ����-@�W�V�_
]���ۂ��-Y7=�H>�o�� `�r$�C�{�#��=�on.��L�?l�7���/���F,NI9"]����U��qf�I)�^�.��6f+H��7W89���BFS��8$`�|ѤYGw��N��垁/����&�v�F���#_��4��L�f-����*���������aZ�L}�G牣6�q�"�,˸���7P��&���u�ܚ��Vt�<95%f`@�n<2� ��C	�~WmO��� fڸ�)���:cbA����;��`7��JZ�yi�����CY�Uz0[�dA87�����AQ'j�^�x�k�\k���sU��-��������;�E�,�|bu�2Bꧡ�?Oc��ĥ�>���.E����8t���D�%����:333E���Y��c!ʞ�;n����ʂ���ٕ_S�Hç~Ʋ�pj��c���v�Bρ��B�V����'|�Cr$��Z]���I��L&�k3��CZ�� �&�I$]�$q��.��1�H����p��uE�ƹ������kf'w3���z�:�yؤ����wW�)%��W����F^c��q5�)	spw�*�`���	s�+��w�C:�����7��5��l��0����]h�K�h��2��
��mEB eR�x��	r�zNV����P�H�=��nSs�����Q�c���υb�9�a�m�x�[Zz������K�z�Y�Nn2�S�ꢡ���u/��g��Q����[v�(b�:X�����(%�@�g����J ��է2UU�ͭ���دe���_88��ýR����5מ�<9`	��t~����vo%�tծ�·#����Ė��h�?����*x�,Ql����n�1]���Pʍ��ׇS;�՞�-W�~��QG�>c�	xw,����W�+j�ZZ�N�Z�����������Eq:�)�]�C���^>[�����d�&QC���-oQo�7R������x�4����	�L���2��X��6\EE�Χ���_��l�K�Wy�^회�� ��W���Y��=lU�[O-5��켹]DCC�OL�J�T��������_^^***~����%�K�&���>24��i4�����U���N$�:0�[����h�~�<]��H:&?��<�����G��s8/��ִ���NT�#�#��kj%o,�*����!%���6.܏���k����y�9�;��$�D���J`_]�3�W���$�L�IF�R���)�M����R��ks�R)����A��]�0�fԲ#:=�[��"����S���E9�K3��J������Kw|fm�΁�m���HYY~GGG��S��1ii�jjj�6�����h5��{}�Y�r^>:RL
��\���Q����$�tm}g����0N�~�/�
��/+�hõw���y���X�)484�x�N�h���s��楝e�J�K;�~��n%����Z��(�ؒ5���q>��m:`�8)dr�����Rx�sD�d�#~֤8-�k�N��)(;��E�"/4�U�Lѥo[���t�J�KЌھm�3�̥��,W��F�o���s���uuI��C�����E���_��,h���V�D�X޽v1�l�O7���z^�9���h��/,LBq�K�9�)�Xy���d^%41�آ-�����3����/���(�E��^ǝwp]����@�&g�c�@��p���.���?*�:[.��R��Gp����	Z8�jx��C242�/ Xg�hk��[���l�\�ÝJ��X���-Dp�?F��z<(1�2��Ð|ˮ,Ža�1������c8�uXU�ta(��n%o�y�}f��_GF>�,7O�[�@c$,�:�����p,�VO�$��I��L͋j5�ȢER�}���Q]�.�R�~�(���Ypv	�X��{Y�,�]"%\1X�x"�V2ڜ�QJ����\��p�n���::���~ &!����N?88@si,*��_��إ�C&��|0�l#����wG�#�!�Y�.UQ=���!�܍�����D��f�%Ov[i�p�8�{ �x+��@>�@����.a�(%�a��1Ypo9��[���{��-��]��~�zP>�������C���Ȣ�)'�JKU��۟�S�cI�F�[n�)II_��f���2�_$�F��a�������IJ��R4��$����l��R��M���v[�.˶�,�|=M��K�ĞE2�K������y��P����~-��"� �#P���E0��� �㡍���́��������u�#Vθ���繹9J]���*Áu�KĶ�EE/P��bF�`h��<ʫ�W��B��J��v?1���vB�t~���Ng	�@~Wq���劣���|8|���F+�F����,+�����]HKKC����|�E����_w*��|��o�<���rk��$D긶
�ѽ3a��N��A}��<J)8 �Ƨ�iw��.k�%w/E�35=�-��������%l���a��-K��,&:�1M,��z"���J�A9��9�N�"�QK^L���{�/����:���}|�kW���\D�F\��,����`N]��4h��KJ���Z׫'PIF��<=T@0W���!��)p��|�3��M߯���% ��G��*z�$a��,I�TNN���r����6}��*)��^�6ͽi�����y����W4���4�o�[ʀ7�2-D��g���4�J��Cǣ�!Ux:�%��F5B��h������w#:4|��Fw"d3�Z{f8�S�	�6g郼�=*4ͅ�Pg~*W�l*��cI+WuΡ�h�?)��{�`93/7�~;���`5{ƕ�	{ccj���B�,(��5�t��poH��
) 6%��=vihj6~R�N�xP�Za<"O�O��l"P���LLL< ?�e�����jkk�¼��"#'7�"�h�(����}c��!.��^�y�*�
��򪚔���wn�jr��@Q3�*4�m;�K��fw��64�l��H�'w_
�z��f&�B~�K ��_,L	j�#7�*A|v��z@�7�#7}��-��J��IO�/ߩ���DS���]��܌XmlX�<�-,���T�����T'oG��+�wխ�kl�<��ak����\I�[�� ʞ��F�����v���V�;w����}�1�54���_NM�b9�3D���p)C,�]��7��(�c[_��(.U67�m�񕎛���.;%	󨫺?=�D%ŏ��<���b�tb�u�C��!L=悗]�Ɛy;�Ӏ� ��Y���ı�����FCC��2(��d\��ʓ1����f_7s���'���6�N%T��H�'��$P��L�SP7-)	����0�!�muY�P_� �(À����aٯ�*��3�I�����$��X-ݟJs�����%}y���Pl#]����H�^��lh�CKV\c�gFz)Xmtv�� ��_
Z�Q���SS&$��	P���9����q�޿ѻk�3iƦy��O;PVm"�V�0t�4�"c��vb6>�S�fO��OH���}A�NNNܨ���66p�a>5x�?�+G*�㔂TXob؅!3���~��J�V�p���t]�fL��M�^�si	�7/OIM���#��e7�NS�|�#�68j���e�{�G�)|�hY�&�27�9�-�����xy��e�J�d���=�,�qVw���Zb]�~���Zd���K�5�׈ή��}�[v#�@Vh�ߺ ��*}��jIy��\� ���ͻk�q��k�p#yw&v��G�=�&]Ue��������Q�����H�������Nw �X/�T 0��[�3�O0N��A�Kt��nta�{��hH��a�>CWJH�q��î���[��?:����+����� �ʴ�g���o���u`0EF���8�S����[�Y�R���[&	��]�6��ArT��� �G\R�.T ȫ��Gھ�{�;�.m8�&����"��k��B��i~�^�G��G�.+���'-��A���;�8}$��9��Ai���:�T��9������7�բ�^^�����,��됽,��h����k�_+lX�F�dNƂS���ư�LOL�#Va ȜMJ�ro\�]i�W�	.���\	�Ku�~�;��k ���X�R�e��X�R��*�ܯ@L���;�����ϗ��ccc�% @�Y�����¡i�k͝����DY��qI��L������G���f��&<Ŝ�����zn��]�F��%�X\0g�X\Ԏ�����X�#����r��y-�j;S�nɿ���i6���QÝP\gM�]?6�e/���.p'�B�Ss�G��)����h�<�����i��H7��3�$�l� n�ŋ׌�Hu���n9��Q>*$6�gƮ�KOz~M��	�����j�]5�f�GT_�梓�Yk���o�(L�����p@1H+"�������F��ӷkh��]&�\ڦڐ�Tv��+�2B�) ��j�D'�T��)�e�TN|LLLGG�׋ˋ�r�����@����u��y���ٛ��b850���Po�ހ�K8��Z0���b�ā���n�3��(�K�N�s��M�pr�8b��Em�á�G/��`�oMh���G��Ud��(cb"�e�w���D$e���px.a�|Vt��Y�[^QX�S�"�X���8�JQ�}�Տ1f߹w(i���D��!d����U#˗�m {l����U���9�/�#���M���|3x-�~>u-��[`ڕV�N�����T�;4��\�d#0�_i�!Ub��cS�1��mhFI�To*�G�d�r�k��t���;zM磼����x���T�B���:���"a��t�������٭�4���M��i����]��_����iW���t's�&�PM�L�a���U����Hv���t�=���Z�RR~gˊ�{�g��~�:��w�?����'E mV$WVy�"!�sΙQ%�?��������BcHM�l%>��U�Ϥ�C֒ 6d�eJ8eb�
k�E}�G`X�^�Ά�c�� ?���Zn���;)��
�#%�ņ���(�����A"e��i���9�:S(��([�~b�����;3�o��q{WD��fx,�����q���������oM�U�\+�8R<��Zv/FM~��PR��:l��S/���U8��ǔ�B���Ѱ����Nk#-:<�У�q��lE�=��ʕ��-�ڥ� B�bs��h�㋵j��aR����K�ei�ZX��������_��2��I�[�E�h��O/m���/��@~��NK���.�υ�^v�FO��6ޞ�?؝��*�_��y�2/�s�L %�_�%�x�0�.�0!-�IM�R=������5��I�vW�'~�a�����D�!�����D�Ѵ ��a�h�c���{Ly��o�W6qP�F6��3�8&�Z�Rr=���"0M������^vW�{��Ҩ���2�T_׬���d�M��{����"PUU ]m�i
$�ɯ�7��a����Ym,+��뱨EY�VC�A`&�_���Z4lD=I?�� 78�F}TU�|��)F�-��(x��k4��"u.�	��h��Y�~s����"�5��s5O[`�F1���i�b���Y�a+�Y�?:�7��]\�ul�mj�	���4Um)�\�HU�:��),@����((H�<߆EEr���rlt;o덙��V��-�R5 ��U�w$�~���'6zФ.C�����p@��;ۢ)���d5T�	l�F�	ܥ�A�D�#%D55�Ҹm�� GK͍��ZN��W�dY�s���?To� ����興��t޸�&>--� /AZZ?�Fo��D�u������Q܎U�A��oџjs0�Z�|L��'DY��c�.�����FC���V�2`Sl���_��q5�E�|�:é�W��4���s��P����>��޶
F7v�W�֗�ư�����n�;�6V�d`Cgh#޳�ϛc&�L��!<d�s9�pر�qn�GE����r���X}yY� Sl{~<�qw47cO>��̇�\k�eb϶hB����	�������1/^]���r\!/z]������B�������EE/��Nb);?4��Z�T?>)�,���.Y��ρ���7�.� /�κ�ǐ�"Ťr� �Qs��J�ȑ�'����;��5�����S�Kѧҷ>�Ư������ʃ��� =��EO�k��|c����c�#�jVuK7���jk-p\�C�����
�m�����z�\�oN�#I���L�3kѶ�-rL�����l�o���/��\_���x��Z4nD9����a�Z~B��_�d�l͛[���-(��>?�ڱ�}`�Xȹ->70<xu-��T�-�*R�)���4���*�#������%4��P��U�4��#�	p��OJ�ys�������Z\��lDdXB�T����c�������jɹE���G%�͠�<5|#!�N���D :�
i��e�ZrL�Z�z�>�f����m�zN*L�mf��L�Mxd��]�����q��sI��:[#�0o%�,3�̋/Б}'��J����VC'B}xN��R�zz}!��d���<㳜%��n�s���i�#u����G�w:@
:�f�����5㢢	6��g�����#��Cɽn��Ϳ���E0z����]ލ�]`��N���皹#�;��}BR!fy�+�^?��f���l�2y�̘�eݓъ���)����|y�<'kT~�!�Mo�X'#���,>�x����?���!��gʹOYzh�.�S���	�rrjy�ʲ%��/9�Z.�X�x����M�ܸ�D}Zųa;e3�ZN弢��$��Z��s�-o�ef�[㮲�P�:[����Yn��n��{��9nᲮ�:���:zɫ\��?6J�e03��d&t~>�@/<�s0�}��a�ƺS�Xa��D���9��%����C5����_H'!��l�������,��/=&~
����f;9y�2���e����X�XI��ᓇ/�Wv;�IyǍ��|��ǿ�!�r��#���$n;i�5�fD�-l� ��sY6����%����g��
j�p:X*�x�7Ш���s�h[��VU��H�A���%�������lf�Ui��^ʌ��k�0�Z��8i�qfeu4yNP־%��X�G������V}W��㳓yI�ƭ��P\���n��ƈk���]u��
�#tF�󸱗�/ݝ�X��Kf����E��<14�	��"��ϰm��;Ty��MNA4��O`��pi%X��=�MZ^�N�`N�j�\��T=(?�����P�q��/2�b�+��xu��B}���	���F����l�l�yT`��#G�e��{0|�o?�a��-z�Π�8Z2���FN��ELFo��s�?C��{���f��Hn���P�
G_J�i��;xHg�͙QK��ǥ0�c���b���dj5�*����N[���˒V��0�ABK7���-��#���e�:�W���)*g�ȓ<?�V���y��]��k�f���ȣ�6o��s�g�_��T���B�7k�*���D��=���򠇌�'���#$7>��������$�c��nr��8��!��tv����*�FC����Yz�Ї �����bE�8��Q4�!��l�z};Y�\����uY�Do#�i`�IM9.[x��}�{�.��w~�׫`A9T��Q�Bh����<���G3?2�n��琗C%���u~b/`sOLLs��wޠi�S']�u/M��ƚ�9=�shS�����]�K���ɫ��u��<)��m��= ���濟m)B��5��9f��x�[P`e2�<�%�QU�p3aْL�`�A���F��x�3�>��i�V���2�?�~�
����Z?��]��l}��L�4�6�%}l̐�GL�*���{ֱq᪫߼}���N=��K�'�2B�b��%�b��o�ӿf���S���fJ�+�Aϴ��u�J�nnBgg-soCB���n O�i�ge��P�[�X����H�&[+5�^����	�XR���S�\j�9jU��<�pL�O��{4J1��fAP�ɐ 9y=A9U/R�{�t&��+���M����|�a�O$�(�N�d�2�[x������;t=iR�XĚ���8<�fw�@�TU�~��Bw9v^]�cK(~��l|'���F�M�_�r����9�L�qP�`���������b/ M���E�c�~��!t�٫�gF�����Ü�#����'A_�:��YQJX�Ŋ�fNZ�ë^��76D�`̜��1��Հ`lp�z�. �7�8F��N��ޓ�n�w�{�d�H����r�o�+?�M������(����r���������{��gV����IPY��-����e��D����lQ��E���.��M��jF���m��%�P��l�������)���o���?�S�G����rjBU��i�����ʬ�zΗ�[�_dTF=�~��ܧ�|h��=���_p�~�S��KHrllJԀ��������(�S��PRNh4xO�����}g�Ҡ(�}|K����#�A�S��bSx0��M���4M�[��\$mmB-ddQ�N|����nW�Mn�E��)	7��'�g���72��Д��������#c��9���|q.)y�뉚�G������k{�mW}3?��Z/+ꚜ����� Ƽ+a�G�q�ҬK��!ź�}��J1���_��>�--��|:̪;�h��	��|'AS~�#wU�o�Sg5�������YP"Qt��p�N�o���0#��}�o�#00��M#$<g뭺�쨢t��.zKu�i��%���8�r/��ZiJh�y�?���II��g�>>v��qs<�V�>?�xt�� ��]����vcf��Z�
�H�ͻ<j��:�����6�>�OTsYԑ�3�B���81@o��˙������VK�Ӿ�C�O��<_����}��,+OuBw��&�|o}��4J��x	���5	Z?!a��q�	Vky�Dw�����Q4ФI���(�E�9B�\�t˭��q;x�{9�|7���R\�f�b�]p�ǱxR���F��?�ء�ў�����<�w�Mq9�u�z��Y� �ߝf�ccJ��, ���Z<����*,�	�(gt�οH��s�v_GJ�T��tN�����.�LBH���/r۴�xϷ�wH����D���gT�_q�c��[M�7�|��9̡�d��^�Y��=�>�n6-~V��|�>����}�K��}��,}hY�V���J��|�@/,6���v���v�|���?��L�� ��c��}��D,@� �P�0��Ě����]� s�^�d=�u���|b͐#���#@�߬�ɳK?�G��hy��z\�kU�	�߲�z\X	y�HJ��Zp|��hy8������Tc��}��ƅ{�
���N]�[��K���&����|K���+��E��q�VV��=�@��C!���vkd>S֫�&q�P�)� ���B<�ץ[��j��p��6�j�Rj�-5ZA�Ңh�ګ���ޣR*Ek�*jS{Fc�ڛ�Y�X;���w��u�s���s?�����rCOT�����d�/y"�w�a�,�=o�xL��ԍ�5������L!\�He��n�.�b̰�-��]�����pm�������/e��)O���!��/-P�W1S�U�n� ՠC�i6�����TX�F;��r��M�DE��:�>��jFh���4M-*�R>@�^��7=��h��/	�Nq{
9ص�m=V���u{�ty�bE�_$h$��T1��`�S݈ۖ�$NMϭ5>����M�NPlE]
��|@�K���b�>�����v�:v��kI ���.�}�=aZ\H�	�c}�H;/H����
=e/z���;a��S+�t��+ɥ���%%�ŝ��['M��l{���%z8��1U�&���������D����O�U�u����t{�箂�(G�a�})�G<)m5#�l�f�g�{���������~��Ӌ���Թ����<���L;����%9g�A��ASdn�u��ww	���u�nmL`E?� j/�T\ؤU1P,��W���Fs��o��@R����|�3ϗAǊ�..p�X�w
T������+���ag�A����i����u��mD�J���M���>�Fynsm���������������(#�6�57=w�ƛ{R�|��j��Ȫ3肁�yn$���>��5��<�:���2��;��XhZ��[��=$�3v���d��GOAh��3��H:���`��Gl~��0�l3+�%�� �"�ߥ�&I�跻�I�Bl����1G���aJO�j��5�T���p9�6�_�����;d��.D�l��*�A�ǆ�&te�����I�~d�S��|;|�j�>���Y���aYX�l��|9��BS�
�_7�^tpf�M��W��2	����@`WT�y��@�i�ڻ�%H�1:��dN�J���
QE����z[����Q"�J��ަ/�n�>�#|4���)mC9�l�0��}��~����iy*�r�qr�X���Ow�=BL�,�Äi◂�<kQ����
�.\� ,IJ��Ǉ�,�����G;��a���FE����R��n	�.�|~��ٺ��mZ�z�;>�����n�51��ދ$/�, ��}M��z�NmYw�P�s��e�[�?��[������9�?4����~{s2)b��d��q��r�Q1�iWZ��/�'�{����0�9��h.��6��ϲ+2t{�u�$e@��OI�j�V��i�"�A��R��ޏ�tK� j��Ek�Bۏ����7_[��cϚ^�ۼ@Mv��Uc�r�.c��*ۂ�ґ��<m���^)a�ׅ�������'_�d}�=��z�<�Z�
<C�]v��_=�l�U�.��a�������֋�j�	ȤSG���ZN����+dW_��+��n��̡��S�8�sk~L�l9/�Q�q���?��R��Ez34&v�����s�K�m�(V�/�N�	�H6��w*�@�ne㈥��"ꃑ�aۋv��K����\%ݠ�S��NdX�N��B�˻�6󭇒�a��KR��7[(�/�7�p���'�X�PQsb�>�1MـF�@U��w�T���$=��,���o�� �у��W'&��(��ƚǍrssw7����O2��'o[0�e�ff�N-��,֯f,M�@�{#��Mo���sAh�Z�mwv��V9]hF�E�(�m����;l�oߍ`�<�連!\�卼�����8&ԑH�,�{y�I�_�Ī6��<c�=�b37&�x�-+ߴcB�~OZ22ڸ(�Ƴ�JA�c$Dk��u~��l���jBo�B�f<3A�����9�7�ݞ�	/փՁU����Tһ�"����U�*��{��{�V#��/?�]6Kj�aT�'A��Qe�vttt���z[��:H��.7�)�LB�ol�J�.�K��J��x�3Q�zlW󻺓>�9:Z�?Ueg��x��J6�FcO����_��ެ+�4'{U���Ur,��49_.z��H�w�@���k��<(�BΟ��~����[����B]�$�Q���[x2TȢ��=$��x!��b�z���ť���� ��!��8�/1�O(<}Wӽ��"~���V��F��<Ks�GGO��{�TG�|���0�4¶�c��}5�w�Iˈ��1#���杬�1�����H��͝m#��uƚ�wwd�������Ri
�hɔg�z#����ygGO��`�a(��0����?����t���CO��˽�]a9-�g��>i?w�����ܜ04��ּ�5�U��߭��}@�[��NT�k� �j�J�v��aAry��-pt�o���t_jju#��j?�V�н$��a��&&�Uzr�d翚��.�35a}0Q�wb��z���^��S����!��-I�9����o�;��_��&$���d��3����� ��=9W�6[��}�@t�#�.zͰ�7A�I�}����tkҖL����^�\U�v���zHPv���t��C_�6��/���1��(|N��Y�tKn_*�+_���}j�Uڀ��}�'߿s�D��a�r��v(�첟
kgm1R���_z:�)�� ��n�)g޲����_�S6e���s��k�Aॴì�=��qt�(w2?�����H�p#*��ﳁ9��'����D^#q�ûNZQ�e;C�࿙qm���e��vGߓ�O�VV��~�s�O?���L��>8���HP�ʞ����{�F���7������"ka��t�9)���jukb>Y�7@j��~�&�Lt���s��+��/d~�	r=o%�=A�H>�u3�
��0�-ĵ�Y��v([+�`�<��Ρ�r� �+�7E��K��#�y�t�>�-'7`S0�3���_���q��{l����H﷾��.f#D�9��][��'���G��ݧAS��̲��V�z� 6r}� �Y�UV��:�ft�Ek�ũ����dK 0I��r��f c�������ި�f+5M�������H�G��s�ϗ.��$%B�H�Z�iJ%�~)k
�����ijz����;X�.�|Y'�׿�K�s��F*5Ȓ�]2Z1� �q���.���D�f�\��6�q>���X��E���ѧغ�(=Yݛ0�����|6F}6�]����)3��t�����'�<���W��l��$��Gߠ`
OKcٚ���*��X�_�ׯ��Ϸ��m� �kgo߼1���������eI����|�s���\�֟?��eSY��#�)T�[���7�~gG�����C���ۡL�'��T�d��5�Q������I8�,t����������;[\�S��$����f:;e>���� ����] ꞈ�O�[��~�󃧶���sAs�A?OV�JgM1��%�=@4ңrn�.ηI����"�RH�{�������i�k��Vp�Ki����\i���(�r�뭩��	<�}y�h�2������X���Y�v����":,�RD��O��{�p����z��E�
x �l�g饮�TIL��	�(8�{D���u@7^]%?%x�o���y2ږg ��ϟ���ud^ڧr�$��<Y��>`6`�1�#_�[��U�_�6����R��n	�!���4��B��1���8���ruu���	����o�g���)��QO	�ذE����xA)��x�ߧ.��WRR���
=�,��c�;���M�V��v�ZUV�#j���f��z�f�:h�	��?���[,0�&��>���- [���x}�w�������`�u9���<���+F���e+c�r�|�\��[DJȄǑ�AG�4�x��k��J���%T#�����\��x>>>�Ϟ���]�'�z{��L�
���]���+����{�z�(� �d�  ~ww��*�ܲ��7E$ǠU#U�bg���O籒�mЛ��РY����{�o�#8��3O��8��~3�����'F�f6bt�P��	�U�5|u�n`6�!��5��ej��j�$������]8����ew�c�{��L]i&�S�``�a���%Cϯ�ၱOi�P�ؚ*x�2S0��\ʮ����~2�S�Ć�~�\MM��0��O��\��c��v�kSS����;��t[q'B>ؚmf�GR9������_��t���~o�6���N��M�6<��O�2�џ��-�Qm����6�I����{W,��9
��;:�E
�vBd��3�����F����q��%���s�ak���'5��PZ�H4/�����+ʙ�_T�����ݴ��)�Y�Qh]݅o:h�C�}9� ��XIիD|���0+E�gT�x�H_O�׽�Ի��m��ܑ7e�}ne/!g<:�������Q��X<��}o��g?��7<�g1y�yx{�����wѴ[�i͍�i3�&���؍�\�| ���FO��z��)���gņ�;�E*
b���^Y����'�C'Z�RP?#~�����m]��X#��w�7��7���|�'�?z�w7ib?�]��P4��W�s_��������E�35]?@.R��"[�^`�A�&��cX��@�ΉF�b�6�W�Ձ/ؠB%(l�y����ys�[�y�H��/S�\O،�E$*���-���m�����2�NW�'��JP�����I�@o��.�W���|�z��ml[���۽e��U����)���P����Ǐ-��^.�@���>�͘ꄯ�6k-';�¿zlj��=�n��b�5e�'+4�G;^�9�E��ux�(�S��3?���'�%�A�����%��#xf�A�p_�)no��)�@���$��t��@�LU�������������Ҥkyhwx\�J��j��N��)���*st^r7��N,��༡)������׽����ȯ��ŕ��:���E��rgˎm}$�eߨ�d�r���9�
�-S�p{f���6�7Q#��se�3�!C8㘖-pj���2G����P�W9�B�������^Q����{�y��+`/��Ɣ��зF������ʐ7r;��<�>PJ�2�
��Vx�V������J�i��h��/~��MW�������U�?�3�m�Q�A�D/�YTy���ȕ�bA�
�P^��L��ɄdJ��%0��L��P��uS�W�Yr�z�������"��!�~�'� ���4@	���ʹ�ݦmȄ���k���'�ki ���y����
�ѷ�35R�5R�ec�4�ö�'+����<0�V���e����SdsT��[)U��+����˘�9��A=
t|�,�sE=���_���u��p�۱2gC�͗��bU@/'oּ�c���Ӊ+��e)�	F�6�$�O�WI2y�n��I� ��R��p����A�|X�P�:+�����M>o��nպ�N�d��_���-X���d�z\В:�=x�f����Pbyua�f��;1�e���pG,�;����\�T���iv�~E% �����wdv�?&��&���`��:��������3A��B���̱jÞ��#�7䉕&�z|J^���n��U���O��L���3��
����G(~Ю�dTZ�P#	7�h*��bNwZ��2��(a�`f)��>Bu�{�p.^����B�ѱ��a�;��p`z�=�0y��>>�8Vʵ�c�:���i�DrZ8?$���+>���5���JR��ڞ�I8�m������nz�DӶ���r�8֑g��o����1~�<�E�oR�G:t�Ÿf�ԫ� (�E��;��w�Ʀ4¬+��Mc	�%�.�^��<�@�jͫ5���|���_C7��<%��9L��t �#7jj#�
��t����_����_l����39Q@���S#x�� �Q�Ma��s~B���j�F9��ɜҾ���&���m[1oiD��G#��Jv�dƔ���"o��!yML�>�@V�֒�\?/���y��6^u�#�������n�������Ѥ�r��K�;(���xn�X:��+G�z����f�3s���cc0�%��ׁ�1x�.�����GDu��RRXL�S���d.n�j���
i/��n��6S��]�2�v~
�O�E�E�r<��e�_�Q݁^'HQ�����ќ�
�kh��53�� +T�|f�4�!��2��P�oB��>✘x,�a��e���#c4z�L�dH5�±���MN��o_z������Z���=��%.z�U���5/%-O�����RB��6�C?���o1�4�"Kb�Q�	���ˍ�ל�7by�S��R���P��^�~��kV�|0ܢ�!A2c8��֧���V�G_��#���  �
�X�8WHH�h�`�����^\��cRb�AsSM�P�"����ϟ��0��������g;G^P�{ J�%]�&�t����z���}�M<?m�� ��Tp}0γq��ĝ����]�#c\��s�����MF��Z�)|���?c��h�����jQ�w�3`V.��%�{��2c��,�,f���K@ۏM�N��u�z��Cl�4���_&��3�m܍��"�,��(\]��ѫ��ep#J����zTo����tʥ�q�{(����[�lv����S�=��Θ�����dH��A��²Dz�բ����TZa���*H���VDD�,_#��.oT�=�2�����?i2�3?���
T��DY;���cD�Jjn�����>��XZ[ C(��z�;-��D��o�( ��\�!D����?�7�G$�EfY��N\��H�f]"OR���b=����K�@�O,!T��KGH�AgJ�yJߜـ��1}m�#�3p%Pk>�"$ףP͢NV3�C�g�D�7�[��ĕ%����*VU�ߍ�����7�^�w��>�Kc�$�2��ac�3��!!�ף7�'hʃ)C;Y� lԺO7��n��` <�	��P�1 �,�1��n>�V�~3UؖN�w�~���?^��]�{;9c�`���q�Q[�<�H�$�({&�h������޻�.N��p�z��#�^���M�SΖfоuVu:�7��_X��YgCv*�z<�Pz�W��c�Lx�}��3�w��-�jװ���_�,Q��ƅZv�oCz ��+�<2�x�"��|鲬�-��2��8���mh:�������\#��DS$؁�O+���o(��W��-���kp�L�m��!�Z@a���Ie��k4iR�\���M�?�����5w��^��1�K�-���k�>�^�~%@`/�>�/FR��vDkcf�
.�r���˛�-��n+�wi)��1�R�+��̑le�C�H�=�)Q!�IP�� dt��g����c8	~'
W�86�p�rq]P(X^���_n�q����r�t��w5Z��+����c DU]I���Kj��;��x����[5� �j%/��a�s�����FNʇ]m;ri^�?䋴�Kv�1f�L�C�wzvZ�b^�QU'4	_?&lx�P�ԭ���H�w�Xm��p#Q���$)~�Mh45�rj �Ս�;w��jzS�6�m�Wҡ��i ��$ބ�J����W����}��<exX{~P���9v�~�[���^'�x�>w�O([���ڨV���ъe^Go'VT�����y��F���O	���y�;@��~p�,���;���[=?�q�y*-���]��5�b$e�����Z�%�j��F�(�L��(��2aL���l)+��˒W�:��1�*�ħ����N��l�r��x��WH��%�M��f���A�Q��L��h�eZ+Nۗ�3@� ��Z8�?6�����I��-ҎFQ����vy VR��&�Y � �Y{/;�_�:�D��Y<W��'�s�#<��f-���/�W� ����1����מtV�bJ79�Ke���m��!<�|ׂ��ic�5�)�s�T0\� �H��4D7ܯ�Q�0�����`�x��_ ����\�:�\��k�W*Y����<�9ȟ�J�`��# �x��B�T�<�PK   SH�Xo�>��q  �q  /   images/2cd737db-51bc-41eb-8762-f3273c40eae5.png =@¿�PNG

   IHDR   d   �   J���   	pHYs  �X  �X{�M   tEXtSoftware ezgif.com�óX   5tEXtComment Converted with ezgif.com SVG to PNG converter,)�#  qIDATx���d�u�+wuu���9�LO�   $ DҴ��l�Ғ�//�����o˖,��%�f	H�� #@�<��9��t��s.�}^������*LWx�{O>��+�/�xF�`�5Ci��� ��ɂpE����0�(M� ~>�ؼ�Ϡ��E�h�slyh�lz�k�.����ޏa~?.�7*f$c躴W���8��F����kX'L�{�������������;��|O�ԏ�G��Iy�7�r��f�l�)��ϔ��_��R��zmU���˶ғgsy��YX�&ē�Af\|�j��,������XC�����B����c����
�k߅��,�๸zb$?wD|roS�r�$��%����׭�u���fHL��e>��0�w����q�W'3�����/��'�A�s&)+c1fL�0�y�����xP1�O�^j���-�^�^�1C�ɰ�q���K�pq�mȘ��r�H�z�Ɉ�3��e�:��U/��_R�|U�J��g?ٿT/a�}��=�^�׻�U��;��ں��>����Q8Jl�%���3����9�}`4
�JSN��蜼a&���~���� �qj5Rg𚚘�"dN���T���yo�x@�K�m��~u�fܱ��F�շ��jZj2��.M}�W̐{|���O�aځ��]?����m���w��+������돖s$f�݊P]����=����A�g䷅�Иn/1���V�O��߁�����͙MbN'(ok]g�V!.��%�7���PO99vje��M娭.��T&��&����1_XM��T&�Z�u7��²����Ȍ<��;]�/�^��_��n���y[gF��~��a��g�`�u,�!$��8��b��� �V3b���J�*��ho��4�W��^Ĥ'R ���4�Z�X�U�V�nW9��¸��]�82�dL��Ɂ2G	l6�.�z�Q��.��'W���D0���w�_B���������m��� oc�$�}B'�{��[�j��>���7�N����oe{�!(ťQ��/m�+a�P8_(
���:~9�O����5ÙV�հ�5msAL��KHnv�Q��t�l�� ��UR��1��.�t�Ӭt��V��`8F{U%&� CA_�41,c�g���/�h��"�X��AӮ���E���A%��"�_S>�&u8���ΐ{�k�z�q���i�����-�f�ɑIܮd�_�qkj]��d����"FYi)�������I��9,-�J�8�N�J&10�E8�+��E�(ä���9�X�xnIf�[�a�K����+aK�`���]�h/c:C��L[ZfDf|S�6/�.�������'S��T��<"Ay�����>̏#�b^¼���7C�PL##����`�8�ל�L)�a��d�d��yJV9�������p����_������H0Z�����[�������Zh4/�x�������TF�\r��p�e��lƺ:7�?�+�I=�'��=WE4����ai)�^�xj��e��D2�٫a��ӞP�?>'
��M,a8��A�#�Jǐ�]��8����A�uU��K����ك!�?�(�[��,8�+��8�N��[���Ħ�e�+�2��,��U�eQ�>y�,�͍5x��E�è0����@�W���U.~|c���*�Q���:�M�R^���"C2�)dm�I`6�5Q8��=~�vZ�J�a��#�?�}.4��3i��
Z� ��hi־>Z�E�9�ECi���9�F�/d�k!Ys1�a(� �l�P�L��T\-5�ƹ(��4*��̱83�3?���4e��$�:sB&�@ځ��2�sFe�L��,N�"ڮ�Z�I�.���nRք��8�a��	dсH%����Vem��]�z��M81<Y�3�$���i~���	���xlp>eyݿ���	*��u@�o-��S�#�P����U����ؤO�0���2Md�PVQU}7��~ e�b��Rq\<�.�~S��ȴs�V��*$��]��OO]Ƒ�qaC�5e�p�,�V�,�A3}�@>.ǂ�妭��ýsT�0S���3^�8�������Ճ7.�''/#O�t�.���!l�p#�l�[Mv-ҞLFP���>��z�S+�S�Ȑ�Qgv��(�6�:@���ذ�$�a\�tX�y��'����E�ꮀ�j��3.���|D�������[�aH����7:E� =�DzQ_��1b�9�ڱ�DF�X�8^�Ua��nU�e�HT_ ��U,c^�����(�����dZ9�a�[6���5X��~d2i���V�l��]"�↨�Dj��S�+�4�n�����_�4��f����m];p��	�	t�&#qE����كjFT�m����;wh��xbY��E��*Q_��\ex�^�>7�ya��S�6�`]W��w8J�?��/�]�82��2a��F	J���e���g�+��p5v�� d�zQ�әt��h�%�ؾ]�ӈP(�hTcHYY�_�hjߊ����zTK3����VR.�������.�(�b2��J��s�$��(�?��4�܍߹k��c��b������D�j��� ���h�C1�4Ӑ��(u�p$�Q�ʫܕ�(��Qj[V�y�Qf�b���Q�j���)T��g��t�θ���lu�ԘS�ȋJ0>�*�/.Y�7��ۡ��P�IV��h�L�+/E��G=�~�6��7�T�dX�7�Ջ,�3�7S�E�dõ05x��� >��M�EgS޹2�hքx&��o�����3�΀w!��t^���"��b|��G�P]ی��!�I�ӱX�hѼ�����_oǀ�����:3�ş������_|�nL�cP4-1��x��t2#J��,�d`��sIu�O���Y����2â�-��T0U�`^Q�~������?��K$k��2m�{��a�N7***�����0����d�R�f[���K��8~��X��.Tմ�>?.����e9��@M��><0����(�a������>�?P�Դ�U����R�5)�8}ދP$�&�҄��sJ6�d�(�:'�;�Y"J�_��:0��s�BPD}\Mʛ��ٿ��s�S��B�������h]w;*�u��o�^�Ao��Nq9�1r��I�<8{��ܝD<�DU\}G?$'�/}�&W9��=7(k"%v�����	���,�a�-�9J]��o�5s��S�B|#Ô�+�n�¿Ӵ�Nxb3��i�N���X<m ��/���_�f�_��d���2�_SVz���jS>�7��x83
�i8�er��X�#��I�Y9���4>@�/��0eՏ�,�h��\�_w�6��K���G�����sd����Y���T�[݁���3*O�xLZ)�ц������w�@\��i왨[����ʴ���B	��(5*�9Yۅ�����e�,t
9	��4�9)98��%��d����-x��i7FR�c���|{0ZQ�O�%��y^�d�Z��YA �U�m��o2%�H8Eg���=��Wˋ���-jA�F&٠��dm�|ҫ��Z+�rt��&��{�*%��)�t�?�s3j��sT�����R\q��.%Jq�P��;�2�GQdY+Sf,�1+�������VL��$�v����o߉py���rL�i�J����������[�8��r��|d�|�����&�n[638RjE|F����~�,���\/���%��>����)�rb!N&�^h����>Ҹa���>�jʚ�E��u�ߜ�~w3t�)6�s��
;��nI�&k�B+�[���s;�x��E�$G��\�tg�E�9�Xd�p�k�7�9�:sR�7c�xƦ���C9Y�<t�L��R��4�(TY�m�d�ErzlJnX����vqE�ߧM�¤��_
�CjcU��?��)�Z��F���9e8��I&����7"�Ί��O�4d���$�6%�ϔ����	�OŲ����+&q�ÏjG�� �Xg�6�$� OZ;�<V�0�̐��Ϣ���6��z�A˖�sX��\������|u�]��_��0'���qiZ��8��'��cq�"�L�T�����PT�}�����1�D-��XY�WN2N�jK���FG��r�:�co�/�k$<��MQ��ϸFqWMk�<��n1{#!�N����~|�ӆ��*rw[=�{�,.M������X��;�� �~�y�zK������oܲ����F����qyҏW����Y&��@����{v������僸��N��85�A��&"1��}�o�/���fū��3.{�V�����\3��V���h���^u��@5�4~��[��v�GQQ�CBJw�{������h�C��]� nq&��/���	���i��۾�D��79�暑)b~d�ZY��~�����=r'��{=~��ױ�wX�m�b8o��R~_�syXf�ya?��7I�W���1���{qcg~���xJ�<�$*����AyΕ�-��/Wҗn؈�/���=nSף�Ģ���ٖ3��W׿��Yy�!���,E�����:�АQ�����f�28��V�d�[8��p�)J��y��$ �ު��CD"��f�Z�vW���Vly
���Z%F1�XC1u��v�W8�~����~���Ͻ�?�м�U�A��P^b������$s	�e���G���W�ƍj�S�Xc�I�RE�l����-Aյ�9vQ�X_
+q�xۋg����Ŕ 6f���5�5�J��+��ɘOo_��)�w�����0Z�|%%�������(--�PJ{�lۋ��!�1$g\�4�*�E1f���uO���Ҳ*T��(3*���+��y�6T)낡���hQ~2O��H�s�"���f5��ֹ%>ƙ��ۋ_�Y+����n���*�'<���5�2591(.�&X�����~�
����qD����FYi7�5���ʛ���j����|�<K���	��*�98Ԕ/U�iH�&�Zy4�L��V�(#*'�[��i&��Ab��E��ň�AQ'��VM����h0*L�\׽f*�?���N1��Мd_��D�~����R>��5�Z-����~"q�,�����*��G�Y��W	�=ј�r��o\]ĕ�����#%�ۧ�j����\������Nq�;�+�k�^;x!��<b� ���w��FD�w���j��!�SJ!�S��&���p�\r��b�0r�8��F���p �̿P�Œ�}]��'�L�;�O�O^: E��2���s*��s��)3����3�"��R���aa�o=��X2�� !#�X陚r;B�c��ӭUZg��/J���~�������ij6]ۂK!~Ef߽�M�	���iF����i=ʕ�ŕ����F�O�r�!<(����F���Sr��Oѽ�>�W��g�TO�����x5� "��`�(k�ܸkj\��{��o�(�$z��#�����"���	qEP��z���^%�cx�L!�c�siǘ�SǑ���Z3��Fÿ�c��C��߾ye����ڎ�^�>�<:�߆R��2��q��k8?>�wc������?c��<���H�qT�[`4[�c�7��kq:^��!j�ݥV{?���I�|�
�y�mE���H��6J���P_%��R�E��ӣ^�I��uI����iҲ)��7u4���J�E��9�X��Z�TsL�����E�N�@V%�I��}�d���^�Ӝ=��(.����Yh?O�=��d	�z�[��'�%�8�<���6Yzz�KKG�2�ej%����Ĳ�P���A�S'���ރ?{�Z}�/n݊�z��]��XU���l�§w����]|lC��q>ea���rO_T&/E�s�{���|nZm\!��1X|'�Do��BAԍ���K9]�ɚfĸf8	���(oG�xnM�C�dM>R|G��4?���Qu#&���o]�v�Pщc ��{{ڕ?��ev�I�$Q��k�'��`��W^;$���߾s��MW��c��i7���tʹ�J-5;�8�k��eD%�0A�8��R p����o��]��z���ӆ���W�ʭĘ[�K'�֮&1>�R��M�P��s�����Y�WOH9�sA7z*�7�7����S����,~A9t�Q"�̸A���UI��Jaڔ����٩^|�|/+����m�老C�4��k���"�K6�:��p�iW��\�N�0���C9��h4gR��aNTR�OVc𬴰H\z���Qlo�뉦0���p���X\|!��_}�Q1|S1�޴	�����ӧ��W�Пb��B���t�)����z��t�*��2٣9��8Y<h�=�[4ZSb���F���/����h`�ɋg�Dw��Dx�| ������и��ƊM2�0]���0=� ������_�}5E''��G��C$�������防×��rv�����CI���58�(�_��w��>�DG�&Եl��dE�;���c2�L4%�󚼤���^F8��)�z� ���&��"����B�]��7���C�B��T��E5{��
e�"U�_�|�I��k�Veб�V��:����]Ės��Do��f��dF�-�O�&�u����=���XQ�Z�6m���'0��⥐V�M��*&�8X�z-g!e1����eI�?�m�]��[׈N�2])}Zd��cJ�3,O���k59�3�&#����5����7���/���^aƎۿ���v�DZ�������a0e�ج{����^�6u�m͍�E�H$��Q�����tm�7���ވ1�@��fl�D,��w��J�+���l��z�2��wN������)�͕I��*�m����������X[�߭�"�=(1FCQԖ;��c���þs�U�C��P�����TJ����醵X۽M��4.'����R�4Xp�vZ��bkV0:epV���nB�)���8hgl^)���Pj���ޡ���,:���[E$/r��Y��>���������Z����YPJ������|��볜��o�$� ��{q��p[������ee9Y%��c�*��
K�%�󘲜��l�PԠ�ݥ%�፼��UWUʿ��*yA1�Wv�Fc�	Ix�p�����7��VL������(���>"����S�L\񅋹�tZ3|�[��Y/��˹�C�tG�vx�.�}������`�
&F.a2�G0kE��{]+�V���a�����lZL��3n�\8�r�ҙ�bJ��Ă��،o+S���ݿN5Y�"a�N:$�&2�7ٰ
���}cH�,�eL:���u"����զ@C�n�	fd�Ǫ�{�N��������^�V�����*�W���ɬ��Š��Mba\�R�3�N�����7 !��:�^R������bV��ad�^J�+�`m�m�P/W>��6x��Mh�ڦĔ�M�Us��>�]T�i�Y�`*����ѳo!���~�t�����C����*1.-ګ�9�yCb����c8�����ء�'���)�c8E�3LQ��h����<?���=�L3;y��V�0�!�vI�O���L\Fe��0蹂��^<�U�����qb"cŭ�Q4�	��i3�\�9��.^�=e9+Mh�9�"�!�U�j�����տ7����\��l�t��X8��0j͞�ՋY�+rU}�.k8e���f)/]4���E��O(��:�� 8;g(WC�_ж���c��C'�F*q(Z�cN�x,7U�=}�	��?`�]�ȟ]��YJ����\�!�+��=��4��X��w���R�%#܎Y%�T���EKQhCX���O��i��.��u�Y�x_ؽAV
����B\����C/��T� 4O���h�Ӝ�N{ m��0�E���.�J�ˌ�	�3��+qE9B�T68�㯝x_��}��-����Eh���G�Lɂ�^�<�BWU%j6�d�"�����i�����n�p�Gz�j��� ��w0��8ӥ�E��sm�m�bE�g�g���I_�KKB1UeNĶ���a�'�W�Њ�Ez��v��+n�U����ӽ�pWJuű�	iN1���1Nhf
!�E� <ӏ�ou,^��� !�i6�5o��H(?�v�B{�^:t5�(�*϶��|[�!y�#b��Sk[i��'�i��б�&ɏPtf3�9�&L���_��I�ŗ0�:c�Ç��jl����؈HD�bd�Yk�n���=�3�r����Şz�rGs��CҴ�8o��������-�MR���֊���d�bc���6�uXR�"���K2��'r��,b����]�ޟ�K%�Y8A��o�;��3�;)3�=���n߈Dx������`$�eh�؂�u7�F�P���T�;D���OC���K��˥�A]�͂��0���Ӳ�J$a�|�� O��f�U �6d
���2��ě������]�]���|�Y�׭�4��C�&�mz��rg�nu�C�c��vIg������qɂ�r���Ȓ�<�9��]�B��`�=��$�&)l��BQϝȸ�VU!�bN%u��*ڱ���^ZC�K�B׮}��pZިt�1�n��5ɰ(�b�7o�,���К?Y*�r�\Y!�&�����7%��X��C�*"�-���C��ݒCg��rǽ��$�2@�bQ6�t�XGt(�}����,��)�3ׯG�R��!TF��RY��i�k�����_gBk@ �Ƽ�@��z�ח�"�P��� �A0�A$G�g�ZC8;�Q�����d� ����a�e0,�(T��7P%f�d�:�d�1rJひy9�2>�OO�j�35I�g�߫VL���@q�ʹ~I�2�lf�~8��׹E���\JWcؖA���6�D���S�b�(	�@]�"j�N[��;�o�,<��1<wb��E��AS�z��:�^\؋S�2��b��h���	�̿|�&��Tc���A,=����<j��H�ܪV_D�����B������!E�>��-x��9��bI�r*\8(J�r��i��+�qbԏP2+zc4�P�c ���}�e2�u�RY�FI��Ա=�R��狪kJW�ҝ��'����cM�w�N'*�|E�׺n�,q:�"v
�ѡ��?��_�T>DDq�D�o�����G��D�	'1|i/����R�Uۘ{��K�����s���B2�ŗ����L��F�P��TΣ?��Иbʬ��Z��U|�y�i1��������q��f\�g� r�R<�Y����JN[�6wwng�Ą��6��O���0)E<*�n��j���ܜGu��S.�JY[g�#MF\
��S)Ԋ���\��J��E���F�m �O���&8�͢�~_ޏ�}V�T��̎���������������P�I����9��:��QD�c-��ڍW/��̌��X�L�V����9��^���������+-xl��D���lbQ�~eĀs>,9(2���wYQ���t��:[���98G��ޅ̒"P:�յ?�aC�#���
��/�)�}<~�$Ք|�=\TFC���PրoxZ���6�_R��"��������U0L��1DS*�*�u�ƜU�/ˬ�� E1e����<���mk��)e���ӂ�λ�51�t;��J�e��Q^�Mq#?��u{O��u�c� U�3rGYu�Dte�u0Y�72��k��g�6�-��$�D<P ���"cJ��`��'˟XֹX��l��
u|�7u��b<`K5��`�&q^&�w�����)	�Lfl˴`[��.�hΈp�
�h���e$��iv�a͔�e�:򕔽��Q��2��t!�b��,e(svA_�LR�$K+��4�b�����QKiC��4��D-���q,w�Vu�f{]����)�({�r��G�asNnOF����=c^|9�|���hɂ�=��dMI�bFYok������~{���옪6^���W8N�l-W>;�|+�K��2exH���C�,�Ȝ�!:��>�L�O�3�ɔN(g�F!+��2HEF\���=W��
�������sq��e-q�7�[�#��ҥV�n�u��h��ԗ9LdK����倧L��1��a����2�D�dRQ�Ux���t��b�m�W��fK�&��1�8��)�E��L��R���3B�E��{�v�b[y��*e�*���rh�c����×�������M�T��hi�(u�Eɮ`m ����OH+v�]��!��Sk:�W+�L�R�{bnN&�G  ��҂�]h/t�f7��U�Õ#�4�嬕���&p�o���+G�1�)~�=���ʱ~���j�fC,��ӯ�y���p19ϦO���B��AX�a�n�)+�
3FKQ/,=��Qq��j!�Eq��:�^T�%�G6��UE���u��s��z,�z�#�q�7[��ժl�ڀu���>>c,�C����P��7�m��h����Ƕ*#���"FUZ�r��vJ)�{���U�Ol��~�X�)��9g�G2���R=��(��zh<�����V�U���uk�N���X|����Z������-[$V��&[����#�+Gwc6����_ ������ �&���x+Z5�-Z�6��в�5��������Z���k�.Jӛ2a$��ݛ���=p�l5���Q��%��KP�&���~�f1�mW���rJG~e��a����yv{#�\-��b�k��g����=un��͛��ы���S����]Ꙕ?���+����]����8�*�*�p��eƬR�.�o4[��=��I�,�b�Ty�~�����ֶ
��3�/�Đ[:�
�ۦ�ei��C�DH�'g�X,���aͦ0�G��Z��5c"
�3�����	\cv���h���h(l�\q�E'��4��R��$:��+%reT��b�7[$�+�My��P]Qt���!_�k�����ա5�O�:�p�[�L�/!��FB@�<3�7I��:5��q<���@L���K)��I1Eo�  ��ҙ����V����Dc�g�W=�U1٬<�d������5�2�l_.����b�I���L֢a`T�q&��9�,$��Br.��d�h�ٞ1���J�psG�o�;�?�����$j:� �S/�hV�'gf�&+�c�,��ݨp*g�l���
I)�=t� �$�ZC��QȦJF7�z�VJ>EY�J�&�N{��u�64��m��14(shp�t�@ ��b���i�6�J'�U�	�T��H<������Ԭ�xl�RXJ�i	��:W?���粪s�&�^���\�S�	ß��n��/U���èm�H/1�9̬W�{H�l�\x C�R��Q�B(9�,:6���)E��B述��.��pK�Q�����XSf��_V�.���L0�+O�f�&�#��Y/ȝ-��$6��)e�D� �a��� Y��[ެ��\,��!���RDLd���x��blԤ������;�+�d;Z���O0�Ƌ�Zt��`>���N���+��{�w�U��*ڷ�,r��W��=�mV�� �.�J�Mf%�|�%���i�(X�u33��B1B4� �/�h�w���d��WYd���Bf��b���#{����DFrKβ�������I"K`�����\ȿ{�0o�6?If�t��z�g�S���JY\�����<�@���ʷr�"E�86�i��~Ά.�������Vt�chS�#��2帐l`��:+�Ӊ��q�I��`x�d�^�թ�,3���o�>aN�Ъ1E�p*�౦�u���hn^�$�q���x�~,���C���G���$HC3+��8w�/SXg���}1���66�*���8L�D�������7��6���5űYD�s�l�Q0����.'����b˼"Kj�a�K/��H��ł�CO�c�ֺ���H���z��ڗ����T���͢T��V���4�
����^�+l��0��"�0�8�79�(wYar�Z���A� W������_�,ZƐf.��c��7�U(�����3��CgD�)�I�z�V�����rnqxQ[����us<V�L�Z�v2M��2«���˩q�qD����$����^��a��t$��LY�W1���a��J�h4��#�)����<�i1�!�>ZE���Q��#=�!�:ϼ��~�J���&��X�IӮ�¡�Щ%�� lo���8�tH9>�c���R�C߆�FҀ�L�pp�_���:��<
gU�����>�9�*����`C1�S��n���g[�|�-�}�e�q�b��o�?5�g��M���[1|r[w��|.�1f'�MY-O䃛S-Ҽ�Ǉu��y�b�G����H��^<X9��5%�q�?AYy�Е��c�]H��\L�q*^>U(Ǳ��GS�:�7�G8,F%YL�ߎw`�ĳx9\�Hƨ����۔�4]��KoD$kn>Ih����[�(�0K	e�_���]j-u:މ�/;���ŭ�V��H�=��b��$Ƶ.��a�=��5�	3_H�n���ـ���1yH�QR�2�P�- ���L�(����i�W��i3�A�P"��@���!�o^\���<�Z]����%���XY��"�2����R[�%�+`�N����1I�V�)��!�҈7ϭ�~p�@1UX�rg�������)�e�]���d�3�5(��8���L�_&VڌT߳���-ܚ�Rf<�(��Z5�E[$XW���h#	����b���4�Mݹq� α��Wvo���������J�Vo�}�a��"����:)�(��+� Բ��<��XDb�RR�غ?����y��������E�X�1��(�yA����`DĐ3�����D=�Fu���rH�ɮ�)�cO{�0����J#����C����+�,W���4T��Y�a��a�a"m�h�I�7i�����MI������S�K��Bk�#����c/�{�G�|Ӏ�ә4z/���Cx=R�X� ����n!pu�]�����3��J�'6
1)�v�℀{Ԭdn��'/���LtwL�*\m���{g�b�0Q,�  N\��7#5�P���йn�˵�	�w.�}�G��n�m.��D�*�n�A-���՝�v�F16ч��������F��P�ݻ'����ː�,���g��	e�P�g��Ր���@�.�UIk�+���UD��9���x�j[o�}��,�m�,�-]MJ�W�J9���>v�m'.)�A=�G�7�~��U4'���8w��;pCď��c�26�5�Bܮ�. �
 ����h�RC���aT߮�j'/EлWF�|�_�-�.�99�(��Wߠ��.1�	~��Z�:��URB�3@��	I���Jq �!���Bk@�g�Z�p�Y�b/̴�)��_��z�J���	��Ё+���͝~�]��J��±�N![��������CP-��s�]/ K��5��e@k̎YM/ւ�W���?�KϜb�}xLT����|�g�nEC���+���#�D�u��N]�Y�1�k��J|Ɠ�$p=��ްH��ݎ��_� q��4���kd�ټ[��߸��
x�bA��1��*�⌭+��! ����g�/�ļ���Bt���dawV2J���+�|����֞��r�U��Gʡ2,�8���#���Z�
�&���tKH�
!O���G�|׋�Nl��}x�ET<�͖�ͥ�X�"�t����f��觑Җ�6� ��պ�!ZY{eǴE�+�~�su�EY���Ν�������_2�q�0��ы�������-�8�S6�Vc e�_��78��u^{S;j�7H���3�}'�/�ꊡb]!2/N���\���>L8U�?y�]T)�7n�"���hFGk���xꩧ099Y�+++�����+�����׊"
���)��a��vE�ֹ�u]Ҳ���]����V��1��Q>���u��X��n��O���k�[7����0��㭈[������Q�a
���~�$�[)�a@�+�a�QS�S�\�R%3Μ9�o|��j������OJ�;�(����$�3�?�Ww��~z����Q�ǽ����(��i�i۶�]ߍ��a,m�p�D۾�'$Oo*������w�\��_������k8s"���O\�������7!7�J������7��p�����<��s���i��� )�ߵkWaW�k_'�A�yOO��_L�Bi��݂��� ⿵�4(f0��O�oS�6�_�^|?դ��z��:���V�ph���^��Z�R�o�iJc"o�^p��޶F`5�E���W�����آ�����?ceLd���������Y�W�փ|���H��z��>�\p�3���P�V#�8:�2�5JK�P�&{����@������g�ޥ�_��}�ӛ6J(��U����B�����Z���L�0�k_�ȼ�T(
_����c����
�4��b��@���MwJ��<+���Z�;4�.��_Af�-2�,�8g�`��}��0k�)�x��#<��GrR��DN�ʏ̤�cu-4�VV�Gd�eMUUUappp�UB��쿦��X��i	V+r����2�|!B��`E m���E�7��ꢕ��{�Tߍ��3�58��ح��{� ���V&������� .���G�l�b4dQ�,+�I؋���s�ќIg�}���Ʊ�v]�O_酻�_����eE�=���۽�J����!8iA����k���'j\k�Q�W����GM"-�˕�w�(��`��x�b���D)��a:�"�1%���hҢ��}��o2�����ۜ�̈́��v��!�1���AF�� |3{���K��|�wbxx?��ϋ�.z�M7݄G}t��^N��9/4a�i��J
���p���#��?���������(�ńcn��&�K�j	�=��+�D��S����T�n:��00&�d���XNށ&_uY��{�l�J��:�b=.��t���/~�6m¾}��U"&-+2Dg�jM�CYc@ 6=���6�/�Î�1���NEc)�r!jq�}�9��T��	wv���c�Z�g��2��fހ�5˝���lڞ�(fL�p�5߬��v�ک^����:Oz3�b��ly*�j���_���w%s��Ї���T��ճ������W@�7/��&q,}p1��\��p)O�"9C!�ϝi��hRΧ�݆b��Fl���G�-1#CY�|�����z�,c-d
V �����癎�.�j�Р3y`؋�}12\�GD��eq�(������~FciX�ׯ�[�����e�{���k�����<tn,��Pl~+IK�-�?�	����!��q���s��;s�Ϯ�Ϧ�!#�j-o/��h������X�$�x2��ϫ�N �\5�+�\�AQUmNcsIPk�)T�m.>�d�r�5�Ϲ��SiFUm�R�lLE��?��p��x0E	K,T�vK�e��P{��J�-&]w;Bx�r�5�p��H.�31��W���fAǘ������Ύ6l�� 셃�Y�x~�^EDY��lP'|hK���D��%��� �~�X�J�V�K�����c�l�|�7��E��>�����˰�8���lW֬IC����𣧺�ozTy�%���j{i�wo��X ��¥d�tԲ-����=tN���{�2�����۰I9�1	�j�KE��	���`ݖ{V��:l7_��~���1�v�:�rYc��e7JJ�H9ȁ����X�ؾm���'o���3e�"�VX���2a\����l�d���g��h���bM��m+��W���_�]U�ƶ-X��^�D��J��,�2�@��k{E&ZJ���FV汶�ag��������s$�m�H���9����r��S�3����)��S�^��}#J�����'t��� e~v[w��t3�����v�~q��m,�a�u���*�&7����G��a�6v�s�A�dLJ�gfO$��5r�#�Q[�1|��Q�ǐ��H4���p.n��.L�hF�6��k9��_�A��q�V��z�uf�'}��l��,Cs�!Tׯ��U��J���*Fч��	����K�İ*q ��г��܉��v�	E�>]|gGF�R�]�����u�q3�DH�_V��?<�ӣ��5���%m��^բ�����Ѳ�6T�DT�Cj���w��ρ�`������n��n�C1ČH<�s3~�kQ'���k���~ǉF{QE<s��:�1:JC�!�L[���6<��/�C8J�Z�0ǁH9�6	��HH�1�I�K�nͨd��()�<�
�K�5�����w������qZ��}2|//Eױ�_���ɒ�j�'#�:�,k�tw�bk�׫~ȼ��Ϩ�#�4B����y�P���K�tȒ�T	�S�n���Z�����c0��x�+�� =ߴ�:/CX}�'=��f�6������Q$n{y�ReW��d%C�+ѧ	c\j����]u�#�Cs
�?0�̸p��/��I�������)�Stڱ^�ڔ���Ѵ��iTd�Dz�w�It�J��,
E=8����I����x��P{$v��!�tf�^�g7���+�<u]��Gz���Ԇ�T������\.IIO�<x7h��z���aei�<s�Z�m�4�j;��F�h>�*j��⫞6x���£g����p�Qb4����uU�����d��L�E�:e��+�V���5�4~���[[�v�G�#C���Qye�\
���q�#�]l��pU��(9U�l��[>�\�	ܗ��?��e&0��ZV��3�ɖ�g�]T��2b�>�#S�zl�z��9X����8<8����詯V4|&���Q�nQ��$���)e���f�Eo)	�	���`V�s�ҎQɶu��g��4e�K�J�s;zP[Q��>���s��>c,�}\'����-є��V�c]]�c]I��w�b+���)"9�����B[�Nly�bHs�ؚXN��h1�����z��3�\n3�a� h,�
�MH���lҷ]�}p��}\�Pu�H����^p_���~TZ�(US�^���ze.�mya/��Ӝ �b��&nB)�Xt��F��2��c���}tk7+�d;;f����K��*!3�+fX&3���L���oՕ��ѮV����DJh�G4�GM�\ e�3V�
P�t��d9v�U��F��e��Ҕ3kfY�>|�(&ٳ��$jc�����L@�j��j���Ud
u(q$�5�
��9�8�؈C��5���^6qX�6�#A��W�/L��?ލ���ׇ�C?F���PQY�A�&b�=���O�P�@g�&��u��A�`�c����^���Ub
�zϟ�"M��[&�1\|�4^�Ԡsb �������y�^\9�*�Nx��g����X��e~=�F8�*]��(Mb����uXj�f'�^���;���6M�:�άNrj3�W�}�S$c��{G��g�zE�8�%�S8w�I_#>�;���O��Z�!��8.3���Eh?/��Hʆ��l��H��k9�9��DʬĒfMh���ݝ��
|�f\�k�St e p�]�RH�P�B6�B����ԗ���x��uY�F��+�`�W�\$�Ơ/�~oH۳o���"3������c���r���n��}U6���T���Pq�u���63�1�)�YՀ$��r�/R��n����F���
b
��}����3E�w����=���=������Ug��f�>V�)z;�}�]�����	q�Ãz[F�;����AUU��`�WOS^��~1C��ߢ���˽�a��mӰcF����������W��']>tt�@]�1{��!��ߋ�	F%����2�D�Q4&,���}����9�~�Lѻ 8	�=��s��{{���p/ܵ�b1z�.c�w�����jf��\NkKb��Ӌ�7<������ΟT�v��qo|C)��"������	�	7�g-����1�f�C�2�"�0��F�6u���Wr��Q�}����U� v��%�����^"\WV�"����$.U޺cf[�n��Mݲ�[$F�P���I��]��.�O�]%����G�/���V�b-ҊbY4f�c�L�m��Ռ���H��ַc�소���5w*4�r*��c��]Uׁ�5۰�wR�Q���Z�pմ���� =��
���*�	�%&T(���dW�)z�_{�����}��)�'|2I��[G�[w�D(�h�EHj5P�:����*��jE���\ e�����f: �t����V�d��W�u�&��ʠ���k�kYJ���},�)��?:~Q�x�R��p�O�Q�J�^H�-
ӛ����Ci;<��о�X,VI�phP���D"_����Vua2���X';~)��3���P�<��K� Lgr��r^�o��
oڌ����o�)�Ks������3R�5H�ݨ�'�Q~�5to�55�i�-�}g0pi�lJ�D�ָC��mM�:ᙖ�I��1CK0��A|า:��GtZZ���Xچ��8ۀ��(uh{{��I\<���{�?�2H�\z�߀ϞQ�\u�h�����˾R�:5hu1��YlM	G�Ɋ�E�Kuf0ӧ?Ňi,��,"S0�H�J��U�d_ĉ:s
�S/"0q	�V�;a�wx|O������^~p0Z!%�7G�hzC+&�b�z�"u�,b�u��Ŋ���|����)�=��� WY}M=��}QN+1Nѭ���l�N���A�@��|T�DZ10�3B'��Ja<k���-�Jʋ-+;h4i9�w���ae�>���y4z��s�11���t�A���e�(����U�<������Y}y��Kv����`�C��FUV��"ӽ}E�}B��E�ď�fdS�w�s3�j攼�c���!leЙ���7�!��U�f)��a�^h=��lX҆Zx(&d�7���|(��3c�b��+�G� P=�ݸ���  n(�������;�[��MӢ�������Tb�r��ʔ����J���0J�9!���!�'c]Zc�=�ϻ��U[����ط"�Ğ��x���K�ja���#���mqUH�;�}ؘ�Bf��/�z��dZ�~��\�נ��S����=��z�׀����l��W3�m؉��?���Bo�:����2Y��Oy�̷��mkĢ f"+�2`�ޒ����)+eFn����D���{�Cx��Ö���kg��l�����x�e��x����h�ޣ�Tg}�0�"(Ґؒ�Ծ��8n��	e���oym�l�@~����bʏ>xLY!3���o�*@��xR@A�����	���s�b�.�b�"d-J��ݬ$� n
��3��۔Ψi��٦�s�hn`U۴���i&��O=��-u�R�I�Bk���W����R>@L)2�^Ō���3�K[�X���D�͊ku�j�z���[��^Bܖ��ʎ��.�RLE�eD�ԇ5ϓ��+�u�w�m�h/�_V1�����1�*���a�\H&���{�}�M�s���܃�z��J��^�@;7W�FÅ���
x���$3�
@ʝM��7��wL���P���D{g�
S��L�r��KW;�����n� �$�g�
j�Mu|a�2ū��-s��+l����'�ҾY��ӆ>߄ )��g5 e�o�Z�"�X[�����T�o��f至��̠� �:�J�d�Ʉ-W�UӅچvT:5h�|΀��s�?����⹊�����j��c?C$8! �&�YjPG.��#�a�nՊ��=}E�M�sc>�2�=�	�_Ly����s���E�|����qSG��rz�'�B�u��߇�c��ҹ2�>�\9��}v�N�ϭ����@�rT��5�����$�S/Ë�VD������.��o�=�]o�\f胢�m	��5ؼd5͌�����&�5�&*�F�N'���Q7�F\�#9�J�Ͱ��N٬�����������h�J��bJ^K\_f��Qס�F��Y4g���xY�n����Wy�y
g�N��^\  ���Xm����y혱����9�T,��~E@��;H�j1�:3c���� �l^�y�㑿>u��k͔9̸~(z}�NI��`) e������4�Ld삊Q
}��Ҷ�˯.Nֵb���2�̔�[u�x!��@�z͆,�Q��]�?����4�\u�[t(�Ao`�q.>��A�V�����c��^�r��KpS���|c� 3z�Q<\9�.W)\�	�x��8����&�xF�!�d�<��oh�Ɔ]�D��^�v��ϼ��3���Vi�b�Hn�F��C�־�Ɠ<�\'fX��y��fIK\�q|x�m�%��Al\�k�܋{��;����Qz�"��i+��Y,���̇�UVl��s��V�5��;>�t2�{��V��ɔPC'��!+��w�I�*x��u�������$�:���R��n Ʋ����a�[>���l�����'���R���F4�-���z�zz[4�c��u;en�Bْ��E���5h�]����1����+����7K���d�O�� �!S�
+e1�\g�a�}Qr�X��ڥT WHc�N-��� Rv���ܱ�_�[�*�ܬ�|�p�j9U����p��  ���[L��R9>4�-M��%����u��]�)י���\���A�I�@k�)��IH;�z:�k�^�0�(��A�E0�Pp�h�d��Q����2��M��>�c��pT�Ο��#� �|\7p̅��~XSm�_4!�V^���!�0!��#�@MC�\�(�#�5
�r��k�L�R�5&'v��T_�o�a�D"���p)nC Ch�,܎������H���1�ܯ���=5[��i+@ʷL)S����4m	�\ӸN�[S�Q���p�1�G�<(�@S�`̉��l�A��{�j*����/��P��l��|Ѹ��L��2|F;��^�)j�����-�]w?������!��kCO��|(Ë�Zt��`�����,?%���g_�O�b�s��Y����Y9���~�r����h �C<�Wr���j�ӓ�K��c ��x߰|ɔ�ĝ�ȗ;�;�"i�-�C�ۗ����4$�Pʆoy[�k��]8�"�B���mx6�,�7���$�e��e���≩�0�q�7�@,k@sIF�����D?��쉬p�o��7:#��a�ro��h�ڬZ�e)}1�n�BkmK�����<��^:�l`U�'�e0?@"����4�>�yL�D9�L�^�D�5�?Ĝ_Ӿ�_�1U���h/����A_�Zl�'g�Oۛ���lnVG3�]=�i5FV�$��U������w�h�9����^=|C�q�)+���ņ�-�,�d
��\ح��.�zx��\�T~v�Y�1@���Jv�R~�Ý{�񦲹U	����aS��ɀ�Ю���_�Y��ϸ��2Y����������4|B��.SJ�Ɍ���5o�PJ���
�8|������R<+��@�,��̠i�Ж5bY�y��Y���c
I#����o�gv�`\9��D��"h6��c�ϟ�'G<�_r���7H�ڲR<����?E�]e)��=�����¿��ݲ��~�Ox����n�G���l>K��cI���	�yT��Ns�W�csi.G�L�qe8�v�Hu�wCx�5�{�S��t�rd���!�:i?����uO�Xb���o���������.�޽Hp1���R�Yf�"K-f1_8{��_�=i8p�r�t�a�����A�L��g�T^r3���}�������g�c��~z�����=x����qebS�2y���t	���s;�_��Ƕ7�n}��&���;��c/�=4"!x]�C�Й۝1l��WP���e(B��^��JW^��MN���F9�;�<�k��.�8tfI�K����V����}xt�Z����⿾�_v��$�'���Aʵ��:��C��b��f�6�Lf�y�"�y�W��uRA��}�y�w�n� ��}�L.yø�9�͵e�q�a�W�5�7����W��A�WNE{9	����Բ5��;J*e!��	�۱�vl�>^g5�ey3LPj��1����YN4��M]�Pb�[����[wsG�݊\!,I��O���Z�+�O�{{�%w�
C��t4�5�O��m�2�o��"���:��^EO�N\���cS�;�3���XB뚏�TMl��+a(��:�5��މ���q<�!����-�p5ʇ����YlMX�,W��e?�@�(������K�{��7�yÄ�����E\ڄ('����ch@Z���b3��x!mWh�� �x<���ާ��-������T�g�WW�Gz�0����_Zp�P1�	J1L����58uɇr%��uT$]u�0V��a���ڒ'R�T*,�I�Y�=���˙�LƑfy��2)nnh����]yp��y��V��iI�۲%���q0`;�i!G���t�L��@�N;�%%L�@��@���f:@&!)�6q�����6�2�й��]+�n����Z����dO�̼��c�����}��}^�H�t��}�,Pm$o~E��%�����*���7�:��^������"H}�]�{��Ú-�<�3�㟞8�}�5���3"��x}��.���n!ru�-��?�S��M�zev�M/�a��k�%j�]8ٺї����Z�i��NV*���Bw�����,�~�v�,�O�[�C����rh�a�������B�V���(�-�<f�&���/�w1BbS[U���a%n}g�(@��e���4ʗ�ӠE ���\��|���B���^v�6"���Q�����+�}>\�{M'ph��~��+�\*��y���[�������b�EJ1�:����,�,ǉ+�
���^β3�Ch��&��ơʾ��*@�r�#r��>8�k�Z�99y�ۑ�a4|�&���B��3C�N�b�9�bܭ8Ϡ[4�j�:�v��݆���p�_�5ř�rn*����ht��f�+6W�bIp]�>�,������g�:<&06A� �ٽ�v�#J�����ӱ���wM�8�Q�U"��xZ��y7�=�l��5܅~{&��\�\�W���#8�Q���B5zcg�ZW�s�z�_��{:���:ԋ6�����;��{���7���w �r�+X��/�`�E�PN0�߆Q�Y��WcLQ�^��Jۧ�Vb�� Vt�W#�s"'G��8�����]����F�����VWh}��m���aDb$#H h\$���AW���i�Є=jq���)�z9zO&k}F��L��v��|ۤ�Π�#�$8ۤ��	vr3�6�)8+g���L�Sv�o�r�U�2��͡B\�R��u�[��}981�R�턅�iο1\,+oeD�"�D��j"<��ن�r�<9.Z�U�HR󍩬�T�9�G8q4��f�>4�S$��b�G�wR���:�o�9��n���q�L4�����H搴�F���H��#GT7�}V �@���k�d
�����Ao�\zT��TK��u�E������T���M��x�����M�[�'UO���Z)��#�S���s~�(�4�>�ͮ�l\6��.�i8�ܨF�9&��=��Ry!5Ւ�Z�=%=^� �)����י�"\���o���<:Yg�>�s���W{���*�2��8�Ӫ2�h?���oFIf���Z��}���`��E��qP5���A,Ms@�a��{0*�(O����E_?nط;�l���-�e��&����kIi�=���"�o�B�G���xщCf�r@���R�0��FM����AeƘ�8��;>����p��k�sE.�D'#
;�{/�\�I�f�%�ıX`wd਌�sԡ&d?�Q(Hs�\��ъlȹ2�jeВ6~��=K�C�}�Eؾs'��b+���L�R���̬l�9�Q,�� ��L�/*4��
��.�2kw� vd��(ï���q�x���x�ָ*w �����kP�|c��F3�\<�U�#�i��\�1nپ6윫))��E�Ox�v���!-��x�	��L�b�֭ؾ}���s ����&��1�q��������yΌ�ЫLی��P5��B7��F��f�ʬ!��Ƕ��nkYی���Q|��[�]����Z�Ҫ�B�M�~�>1�����|����-M������S�`�`�ħ��f�o�EŒ���]�|2z����>��]}ʖֆ���t5o���՚}Y�Kk|����k�j1�G�N0�WqVo��_�1o!|"4��Ng
Y�I�/�.����l$�b4��EK�'�#��k�u�:s��.mt.�Z[S�]�b�,�^Zc�cT��n�YZ�k�]��D��u��/�J]��)��ʠL]'�6'g���f�/-<#��k�n�P��-h��ҌI�2����1� 7�5���ԍ�Y��yvfi5C	 3�6��KFF7��[V�d�²g��Tx��E �eɣa��'1���/n��ӷ݈o���ۚ�:e�-�sm�ǓV�5���Bog�R&�2���NR��v7�w̯ˤ�b���sZ�@�9��U�A�� �%!�3�m���|��'�H�Bn�DB�Dӻ��5P�(3����6��5�*���׭�ҍ��p��24v��V/2c��Ԭ* ^�w�\�ϾHo/z��5:��_wT��n��WX���v�7���Q��z{�ƾg���1��=q�=��Cݓ�B��r��p%� CCC8r��H_h���뮻�m䄑d �� ��7(#���L��*���m�H�� 5B�$�
^��O�ѵ�WlVe����4�?�����IT���������w�Wym����'�۞4+AYn����~]���z����Z���mx������ۃ�JY!{r��46����e��|�ǲ����-����5!#X�k6W���{��U{Y�������D��!x�%t]D~Q��Ɓ���������ٱ��oʏ;'3p���M��K�;aӍs�����ܰ�
?<|R�X�0˩��(��%PQi4Ӊ�0QD�����0�XH0�y�����ڼFӔ ���s(�3j�KOl<׻����[W�Ye�n������fx{y���\݄�SqDL|_��o��sǽ�n�6��Ki�R����*锠�	뤪��>�X� ��6�+��fK�E 9.�z���;�ke�it[�_`��.Բ��i~=��HlRo���r��ru����=��[�7�0�m��|h8�`��H ������2��<I��^�����XV&�J �/�z�E��[�S؍g$a
3)a���H���'�/�s5��ʤ�� ^��!a�]���"��V��
T� �#�z���% ��Du��F�d�&qQW6�K�{�E�₨y:[��3�����B0�z�!�P��� �^FPÞq�k�c[�Pf�
)7�rpz�`Fɒi��j�n-lEma��V��æ�-]㥁2�X���R�}�zT��i���n8E5d�U���3����`6]c����|Q��������VC��G������.���d�>���gݍx��MbrLS{��}RKkl_�v܄�lk�h@L��~���j!3�"���t�_W����;���z����m��ΡT�N�[�@}bX����K�l��:�^��vj�O����!8N��tUn*�C�w`wv֔`��k�������r�U���3ޓ��h�Kg.���R����7C�k�a
It��縃A�	)�Iy�TS�d"Y3��ŀٟۅ+6�f�^���
!B�:��|=������W�{�9aK}�se�v�����`����%�NTTo���C�}=��A�DL����74-�0��Αe����֖�x�=SVV6g�6���������؍�(��`�s�U����>�A���YT,�6��_M�,MG��cˑ.1Y\�l�Ṕ[��O���ە =�Q��z��&պX�YB�ܱc����̍R����?����9�R��"��7��kBc�I�P��|��Չ̴����)�A-�^܁�63�W�HY�7�v2շheR&03�������q�2;�/�\��9s=�DH%�����i$>�cP 3eܖ�p;�V�V�L�-���nF�d�&�O���Jw=�ZΣ��YY��0��wF�����Hvh]\@�Y�s�F�.����R�Ő!LP�%qg��9m�����aY\7��e���E���安"�!ZVk��85Z���2���� ���E��d:���A�#8�хׇ��!хr�z�?�/�r���J�BP�D���k�T��L�����.J���qR���P	V:��v�'��݃��%mm�������[2��)�}�'{���:�d�م�fp���/��]��ﵩ������d�7j\�L� _�J
����Qcb��3�lj���9�<&ˊ�l��T�l2@A����̜��4Y�6`������I�YK�]Q���Ƣ<�ٿ�T��N��_�J��4���������a� t���/Kq�[�2.���;Y��#<���{�~�ӛ0>a�y��Td;�� +\DxAD�Ud���M�R0����ĉ*�w�ܩ�&2��=�v�
�6��� VMM���oM�y� >�����ǯ����:|���زe**� �566��߰aCX{��*ǁ}�9q�]�c���*��[dG$>~*�C��N8��e�S.�&�;�f�G򔘅�i��O:�ʋO�G����ÿ�g�j��OW���E��*�(
%�Ya���>��F�~�i��W��v���Q��3Ϡ��ZG/�O$S�]�jՌ٣�a�����E�����+���{�w�y�>����s����#�<&��3+K�9�
a�3ٰ�<|���^�||8�5�}?`Ǆ��,�>R/��5<������9b���3!(3ΰ�HDr�e��8Z��y��D��bB`Xg����oy-���<�\���^��Au���Α���$\�4����	`#�KKK��k��"	����=/��,�/.AX�Y]eX ��&��`TY�611!p�� $�\�9>9�;�Qc)�uC,D�F�w���E�ji_���ٳ��`�'#�˄	ΐO��g�<#�Ҙ�E�o����E�M��J�S`�8#�/�} �I\"0�^*�====J�� Fsf���ҫ�B���_2'#	B�ub�f&�Է<%�Fi7�G�2��U�q�'�v�?���%��A[HY��#J\��4f�S4L#�+�:ǐ�L�0������o�|�D�قU�`\g		���$��\	b�?��Y���c��O���Q>V�vg7e
q'�G�c��Ĉ��k��i���\\� Dp*�=409�LZ�%�f�7����ރ��@o4DD���y�������+i᧕�G�q�'�C�K΢&Z��O��!̖���AZ�-����px}�}#�]�h�z9�YI'��MZ*��\��1�O�����>ĭ�aB�FsI�U���7<����yi���j!M���u*��E6w���ۤ� �E�Q�e�|�9�V{�!����4Ї"��%p�����1���)0�4�=%��+H�Hgc<0�ԜU���(���Xn�q��v��r�$@�='���H~�+�lND"�'��#o�e~E�-���{�X���؈(q-cL�]��^��Ƅ|��n�M�6�3��X(��+���3����E?��W[[���v�]�vzDOڐШe<�Dc}���oN�(��c��N0� �`�s-,v5�Dx�v���<�܍�[Y�!�hd���y�*q�1G�ƍ��SO���qMΐhGd,0���&Hy?�����~;n������}��:��t�k�g�)-C��M��
��$+fG|~W�s�?�2�"](��D�K��"�"'A��TҀ�}�QC��^Þ={�nݺ0q�	�o)�r~$}��n���ٌ����a����@��ov>�i��'&�ym�jݸΖW_}5&["AȊ�ĸ�٢�]]]��r���+�����L�;v�y6+=��|����('7mX�����Hnmm����!rA�DC5�j,^knn��Ç5J/�n��__�L�M���xg@��|����/��X����=p� �x�pNs/y5��"�Sq��]���E ;�]�w�x��򗿜�pT#4=���g��-W��x����g?�H��U�b�_ ��y~~~~R�׬ĺ�k4Vnf �tP�Z�f��p�'J7����� ��rd߾}ػw�a$�wܡ�Rq����~���l�-�ܢ-:�$\���j�����&OG���O����p�f�\"���/3�J�Kau�e ����$�]�,�^���*�,2H��o]��.���)�xH�X>��]�f�*E�P16�X���C޿"    IEND�B`�PK   SH�X����+  J  /   images/5644ca41-1cf6-484a-bb07-c2f9a6f5b19b.png�WW0 �]-�+D��DM6DKV�Ѣ����Al"�Z���$z����:��V!z�������g�=3w���=�:Z*T��  ����[��E6ٝ�L]�{K@OUco ��� �����|�`>z>k/{ ����x�Z{�xx9��J=  @Sj�r�o3v́�I�L��S�g@`
�\���EG�T<e!�����DʲϘ��|���E-	:3עt�&^7Cx�-��
H%TH��!�U����������C��ח��(���~�|����>��`����e�~�L����E`"#�n�����bng��0�d�w��f��u���R?	X_�B����������`؂v�r��I���ӑ1��ԙ��*3~��_��:a���skZ8��[;��"���� ���p�HZ�������1�d���g/ǚxx���L�	K��%y&�Zt�Q�� PKI�!����O�Z��k�>)�|yX@8ҳ�́ߖ�N��+a�i��?���m�ޢ�[e�O�M�����"si�n�4{f�g��!l�4eqz� 4W �J��(����3=�ͤ�;[AI=�� �Z�G�'�Ci�55���T�eqo�Z�K��T���/���m�p��&�5��(��sց�ѽ��;�:���v��F3��� 氉2��G�;H��1��"�{I6WY�#�JJJZZo����gKJ]����p�Y�*�`��&���i��&�k}pp���F�oʡ�t ���>�x���n�3c�ºk�����Vq�[˛���ai�ɢ�L�7~@�ĩb5�W����`S�O�=�\"�����j��oq[��Z�ޛ��~z�G��/��G��)����Ci�h�k����i{(z��_�zģҕSD�i�����SO���"҉5\�^QY�u��6W-"RoMaJ�`:��󸼝�@�&�GH(��3wkװH<2�wgv�9���>�M(�Ѱܢ�k	u��WKJN>��`�i�꒬����Bfxn'�R��c`P1o�9��T��E̵��h�ޑ�OZO��F~��nL,"�h��UO�����`�}�p�P$v�"%Ʈ�Y7;�>��B��Q�2��'�З��>Q���ߨ�|��>SU &N	�}�C��<&�uDi�ƴ'�5_��i��H��dƱ\�7�[�i�^�6WŊ6G�M*U����o�c|��3��g��4jf4�퀋�Da���B�h�bs�H��Lu���_b}���p��9�ib�h�Hm���I���� ��w~�:�Ǚ��(�Z���iaa��-%�X�0n���4�S�P+ҙ=ߊ����D��BmvI�Mm>���}K��A�U���q���LyKHk&��MjB��}���A�f�)���D}�ü����{����h���xܞJ�tW�&P=�a�kw�m_,#����rׇ�߶<J��V�vg���^���ҵO4 ����l�IGB��L��PS��ڽ�����	�;m�y�}a�.��%\o�jͧ�g�# lF�<���s\RCj�ch.�5O</[ߖR�̔��{o�Zwu��H�UV�E���_�#>��N����1�+��Ġ�E٫�ͺ���vub��Vt���9c�M�j]�򏻏aj�(p$v&�99�r�ئ(��J��Y&躙l��u-�1�}x9��x�=Y��絗�<D���T͢Mxf6���Ȉo�����{�W�������fF��Oʁ�����w�7���C�f�<�{a��ḡ|̴n����*��V̶Q�$��e���YWc8���dO΍��$V� =�z�z��!�Nj��8�H|������~@�����;/4��ʽ}�Btnb��D��WsV�_዁�tPY"ۃ�t�����P��~/�9žcT��bQ�F���n�}kM�F=��(&�����<�{�W���i�1Ӣ3F\QJ�"�i3���%��1�ixjF��aƓ��r�*:H�s�Q�"�@�g�����������$-x��d�۴�D,hO$LDRS{�T����ib�7�G6CK/X���7�ɣ� �)��֚��tWDE��+�9��R�dV\�Ѽ����E���X�;+�[���P�a�Ze�J-s3�~v#sA�;~�sDh	.l�//��ܦ�:�S���Ż��|������ᬹ��FO�����h1 W�f�V��e%����\+C�p��T�8�wʄ1���l�5k�a6�|z��j��������2�zX��:�ϳ9	���P�������@�UlA��0Ԥ����\[j�4�r4�j:UOz����'y)c5�����;�u.S�����t�i��p�*y�0ؾT;bg2015A?�Wj�l��ۢ�$1ye��K�����E�^-����T0���8��� ��p��a
�`h*�Nj`���S�^N���dB�@#�*N�CK����9���R���૕V��v@cy�;�K��z/:�,Xi6S|��궣���M��v]�� &)��\�4���9h����_T����,��u��=�n2�O�R$گ�[?&̽�W���'����>�޸��R��q�ݐsW�t�)���9RqP�`��]�
� }5
B����g	k��g��wf�Hf�1bt��}����8��c�N,���.��)��֩LS ���5���梓EjP�r
|-�������q����F�(���5,�y@� g���Z WMP�;�,8#�]$.%'g�^��!��.�x-z�\��������NQ�{�zAz���Qr�����-wT�1�,T��r��5:}�R��`Ha�ځ_��K��������`��s7}��3���ڑ_�129kzV�0��� ;�#+w7�p�i���L������ xT{�^W(qm���_N@xGY׿�<�F�^�FNz079[WE�D����i5��n����a�Į<�={�ܕ���V�i���ܬ�K��$�GȰ��ץ8IU5�D:9��W�Ռ�,!���%l{)�8Do�P�H�~5(�\@��S�mmu�e�m�ڥs��>+��ڃ	:=s�Cl���Q�X�f	Ǒ�V��a�<Z�5#u&r8▴ ���c����~��?�j����Q�EB���C��C:��h��a��L�І������l�z,.���'1yiV���F?��K��.ϱ����"�lC�&A�{>�v݂���`Ԏ��:���<��Pj(_�q�e�E}��*Sy�ţ��)�E��k�����N>�a��Ȼ�U�Mċys|���_�֕�d�.#pѫ��4d1�&@�h�[�Q�����仚b.��W����M��R�k9�FY=�t�fn<O%����\j�l���t�r+�����Ñ��T�(E�@D�����3jbT��hy��b��A�`j	�\)�v0�	Ăl�r]�_��_�%K��*����d�PS���ſɅ�.��{ӕ�#�X���b�\6��K�g��,id�dQ7�o�|#�p���JN��w��
F�$L���2-x�s��`�
�,"#���ށ��1'Э��x>���
#����-�|a�M��^Zօ�Q����q��>��Ւ����v�Ur ,��[���t���(dN��z*�Vvq��}zR���j�fC�;<he>��4�d�R��f�Jso���|���_����|	.���۷�R1?����#�<=���	�of�d���{�-����k}2`Q�5�����/���q���w���t�B��a�˳� N��%y�{�es!}̰B�crY�	5C���ņ-5+z �!�K��U��9i��hE��������$M:a��Y�UmW���JU������R���)�\�Z�~[O��-#���b���T��\p�������O���h�_�fR��L�����WNs��B����z���{Xc"]���oMe�X-��sī�M�`��E������[���Y�T��0�:������ϟ?�=�
^p�>f��ݚ�4v1>�^���f��"ȴ0��^�f���J�j�M�ZŐS_B�M�/�������c;��[�sCT��#�܆���b���?PK   SH�X��p� �� /   images/7e81f6ad-0912-4ff6-bfc6-e58bb7840941.png�wT���6�qPDG����>� J�@��R�FjpP�A@����& ��&���"=@BB�{��=��������z�g�������>{_��{�s􅞎������@ �ݾ��>���`�t�����1"���mã�8z�9���>�e�@�|�9T��� ����������B��=tu�yd���!��p�8��������_���/"_�c�?Ə�c�?Ə�c�?Ə�c�?���#x��ap3 q�1tS����1~����1~����1~����1~��+���������f~��ռ�䣊ʷ���������N��W�e9��;��Z�����=�����/�̍.����;��'��Xb������jR��Rӭ7�_��tg�WQ��;G�v77�Ҩ#�S�v�P��d�^uw���wE~����1~����1�?��C�qLw��J/i`���[1U��*����hqE��R)Va��jt˗/�,vLe����|�)��*�N}_CW~�����C6om�Iu��Fo]���O���j����Ӄ�adF�� ɜ�)jϣ]�x�A+�n�iz�����T�'3�Ԑ\�c�t5��^�ih�_͔;�o`��&����Y�O������HA2������h�bw�χ��k�N�>aS�淟�~B�Du����X�<�a+l#Z�V��yf�._{|og#����n��Q����:Í[�(1�u����I���7�<�Η}繻���_��ƿ�lB��Qx�ING�^�Q:�`ݦfB���úL�?b>߉g
gVO���$���d�W5�p��s=�[�-��d�z%��`�zd�����S�
�2NU���go���3~ϋ=��#��y�-�-� ߹.�2[��.�u,goz�&
rZ�T��88���<��Z#h_���İ���uX/�sTF�lG�h�[��t�ڈ�i<��3\����e��o0��p{�R���O|��b����t�� Tw���|�e� �')�^��1�"�c�Y<�-a3�ç�fV��A�E@Z^�S^�Aś����-�_�b���a�C�䩡���&�@S=��R`�/n7u*�K�f2����z�̂*UR�Xw����;J���mIW������Nz��p�l�;TmV��Hi��&f�ee�RX�_צx[��6&��4�7k=�k
�P��ah�c�{�h��rvv�����ͩV�K�Ֆ1;W�g���s:�8=oQ>~ؽ�|��["y�8�d��9V���m�T�Y҂�_C0߮mH$�;.J��s'����X�Էe�:Nڥ��R1�?�dV���+'����pזA�G=���3��NP�jc:�����f,� ȳg:<k�\Vj���U�b��h�zE���n�(Ѱ?%eHm$��:i��QyuYK�������hs[�9�v�E�}#��=AYɚͷ�����j6��~����×�j9������%�I�±��Ð�m_X3��٥x�6�4�� �1}*u�:6[ĺ|�i�CI�{K�\��-�ӰO�� }�/}D���d1�6�Ű�Z[��
�}G�2OUg�@�\��n䊳IKA����	��~y��]��>��\7�(�qj�?ޛ&YX���Yf��קּw�r�e*�)��Z��(
|�KI<񓳨�r@]u��5o��
vL_d<�dL�U�և��R����T��@���_��}橒�b::c'h�m%`��t#߿��B2"�'�%��+'���g�ZT�+\�y"j����կ^�ʙ�P����#��{�ld�p1�y�?3��˫.���^+�Zm���u`�a�Z�]��-��]��PA�9�}�z��k��o��ru����i�&=����/(��}���!O�Z	�gg��oQ�7�	�������n#�~1��|ʘ����~7�����V���Ɗ��<yD^��bd=d'�S�$�^L{�ؖ'��1I�v��˯��uYW���Gf�U0"�뱱�u�2�ל�����5��
����j%�7TKj����6+k#��'��{L[~�l�5��	��I��gU;u�,��r�{ ~ G]��$+(Ĕ1�VQW瘋�r5sp�tv�:���n��������%����0�)w9ח�rRRO'�\�|Z�A Ѷ���S1�ڔ��	�@�־Ɉ\]�tV���6��U>�WxG��n�>D�J�9�ݯ &UlX�Ƒd�p�v�a;Vb|�l9aX?,�y =�9\��yI�/��|���Y{ٹK�"��Dٲd>e��k=M2(�R)	�t����A��|��A��msKd�zr�V�@Gk�
�ѐb��m{:q"��s��C�SY�n�U��`aف1ȇ<����Te?K��M�;��Z:�^&��G�/mΑ�s�ܻV�h��{x�}���;�Z�B�~K��ʻ��	)i�������d���:o�~6������s���
���((P�n���ӂ�ac���l`>{�8R��l���+buڶ�j�V�4���9�,�ys�ҋ �R�ᇠQ�.��m��~���ѥ�KYLO �E�<ǧ�RjG��د�_iV���:F��u�[mqkG��N��y�ٷ���	���>~�b�IDW%�*a�$�]<�Iſ"�D\��5m��F̺���n�u�S�I�,�c�U�B?iɇ�	_�'Xơ�O�8Bmx�̧�u�֫��<e[�\��b���|���{�}���>�Xn���E;�Z9&�,͉Ц��]�m�������a�7�خ	�l�"�u��YsHQ'�{g��=��ItouRz��ϝ>��1Tc?d]���zJ�LE�C�}p���X�1�I��.I�J��55Ͱ�lw0�X�Ī��n(RSC��=Y;��ۙ�S�A�C'V��Hl;u�PT%v��١E+X�6�F�H vt���h�I�M\I�&!��/4]ޚ#w��.+2h�(����CV�.�8����s'�k�IY����� `�b�K�)V���UϧJ��_��x �=h�c��&BOqw¶�w��
_!ƨ\����i�X�>�ғ�+�u�׊�wO�y��S~�B��ߦy�9�yI�.�*� ~�x[�(M�����3�����ÿ�󒵔(s���my>��7�C��� vx����բH@ɋ�Q�w�)� ��A��}�Fw�b�+����U�^`au����9GR򘲴K���ŊJ��n��.x6j�����j�s+�g�So\��e��Y�3~S���1+$��j]�����&{hnTM��=��B幖ۗ�k� ���џ=�+�26����2�.�
;�d�S��(a����3���#:�;�K�wJ���Lŕ���Z(�w��Xѕ��a`ZBy&8�v/zB�j��"�i�ig�� �����.��w�eZ33�)hb��< QIi�P49�]<Cq�,��,���x��@�>qJ1�g/�,��zѿ��@奧P�N��*�_Э���ج{m��:H&T�����I2�߾�S=a.�p�tX���S}�]d|�д��P�su�Ǝ?���*({&�w���l�ZHClP��1�S�tMzlMdi6���k��3>��T��Qo�^�D�1��ޠ�~K��]V�w!ҖK�j-ۃ��Ui�뽷��W��_���X�9��0w_��Si���.�s`��Dn]����y�7]̑	��E����
U��>@��9|��7�	��k��s�u����RJ�3> I9;��nށ��0%Y��卤)u���Q]�ޖ�eđ�߳|���bg+��v�O�欪��9�2�� 8��f6!i��}�	���~���VC5U�0T�����+�*t���@�K:xM�bt��ux�lܗ�&BX�ˡ�i�������Hߩ�#�0�FE@vt�:c�dlz��$c�k��2����0��B�m[��:Qy�Hb���V�$�оN��jc�_�0��CB(;~Y�4@��^��ި����>%�S����s��2�ǯ�D!vv��ؐ�1Z^*�!���]�o���z.������M�f>��琾�`x6���o1&�-�;|����?o8r��x2<�c�Y>�9��a��q��T�O�jX������38-�tN�~5M����2O�}�ub��ޖ�0+�����m�uv�l���1��]sT���APH�� d3�D�dQ��^��%g�>e�x"�)�r�b�H�
Y#�"iqYvu��|�����FZ�U\�!=�/`F<��v57/��2�g]��������z��+��&].�p�4e>\�L��`y7��[�!$�,f�k�}=�Ņd=HM9�F��+6��hU��T���A���+���..�����Ld�CjJ����m��Qƿd��2��avj���t|��������XGd��"�[�FN����ؼF6����@�g8$�)��2�����fKU���A�)��q�����$��,�iO@��]��L�\>k�V�Q_t���6d��F~�O��S9�K���& �AR˃�"��S����1�!��S+
v��������6��23|�{Qt�!E�eN������
�{�� �dJ+pȼ
ӛ�������3(?�V^c��s�����n��B`�u��7~S%�Kا�A�+����pp�~[���ԶV�9�~-���
���t�2	��VX�g(�R�M"�?�	@�uGJwK��O��X��YڭU�C �VС0lȖ�B��V�N�f���5�����N�Eë�﯌����������$Ɲ�����
.����^�ŏ�{���I��״e_L���;����Q,�,����8���!��Rkq����Ҫ����m�r���]i/�?C� ���"�x�
�8:ٰ!�!��r� ��_̻��ϊ�cx��)�X���D)�� s�4�X����}�Av��,з��"�7��{�P�oU&�o� ��RQ���|e��\Eo�N#2ԑt��/fӟSJЯb{�¤,�C9p���A|ښ�Q�.U@�;��>�ttl�V"�#6�!%.8-V��@��@��W�����E�V�UM%�Hn3,/=.t�!�����!P��W)C��֍�,p0�b.#��U�l�Ыk}mTz�87�6!�������W���F��BWͅ�r�4��[��Z�sdF�V���IB?�c��`��/��1,WD��')�o���x��7��J�6�;�n%��������!c�5�\�ñ���}<�W�yI"�*B��}����,pl��Ímd�C�S�컶H��z��tG���\��T{`a����ۈ�Pes�i]fS�;Yp���-�/�/~�V��!0Rj�=]P��ҏ�=�|���+B�#��6�s���������/�aH�'ݴ3��@'O	1�\_WV��Em���0�����<���òx6����U��l.���&@�,<�a���=\�Ɇ�	�W�h�&s�@�ջG�#�yow%rE�	']1������E���^q�O	�r-\�;�?��4�� �'��>	F1� �ʓ����jf�9�Ĉ�&G@�Gj��KY��tub��J�N&.��#B��Y��铥fÉ�Tܕ7%Ѡ~ַ�r�9w{�7:�=��Da�WC����[vh۩*�����=����l��V���LʴC-M���xQ�Vj�}M�<�&�C��}�='�KB���q�5[je"F��T=1�ҥ$A��D�߆�6@A1������F�{%2���3j�u�E�Zˊ7��2*�g�v;)_��i�rR�R���R��/�]n=�C+ԖWynU��Q��H����>�=�S)(�ڏ��r������I,���&�(ut������I���q<�Pr�*ЭY�մm?��t�����&�߻�E<j�/�8�o s@[�_D���Ed�����)9\�B?D��V�G�����YU��������%�{�-�R���&��A^�"�-�����X�����5�L0���/@Wh�����T�c�mϰ�+4#�U�����x�`�+���6zH��yaڃ�ZL��%o�<G�;]�?Qam�vg9)�̩��΢�r3��؏0x^���'`�2t���.� �*э�qz^:K,��T�z��	R^��{��oE��}R)eʎ���lL�Z��}��Z�Av�m��^z�,hH�w�]~jv�n��7�TTu㴙�֍5����?�:@&k
$*�#`K[�E�]����H(��@#�J�b#JDNя��8oI���2Y5q�!I�w-�ha�ns�2`N��������Kc2%�p�=Z;��R�\/%E���F��G8�&<'5_�%�ғ1�u76e�� d�!�	3��ų���"Z��X2��`�wfIW� 
Yv�,�
�^���b��X�%-Eos�U�ӹ�vބ��I�A����c Z�?��/��R�7Ǩ���]u����G;J\"�q��_���zǥ����t�2�M�����j�hw�Z��"W%�j�d�L�)��q#�*���gA[��J&ٜ���J�6�W�d@�g'|ͮH�\�{BnC9	��_.�,6�^;��?��Y(	����+U���ŻX{�=ڐq��.�䲷�x.�k�JGb� ���rK�A7ܥ��}�+�� ����#2��������Ak�vf[$q9%�<A�b\:�"<e5���J�������$�(��B�X��Z�JĖ49� �ڃ8�!O��ϵ�&FIb0�-���[�<��n�U�)����y�y"������l[KNEgF>���@t��eT��0n~�����Ģ�zg`KE�@�� ����z�l��o/���=:���4?��Q��st;����m_t���n�/�yP�2���/�o]+�dg�\��X��;�>��$�,��$q9�f�ʩ�R�oA��>�����}�Cg3�0k4r;W���W�T�<!` �r;hv������SP�́p���:��Hն���H�Qg��0���M +n��4w���E>����~i)�(l���T����ڻ�q�M��<����oOOeAC�W��f�)j.Y���b�{��y����<7��6.Wák]b>����of��)����Fa�Q�qګo^�T�JӁ�A�'NT�&���T�"O/hᜧJ��襕���y
B�Z�:$�\F�s�7L�&lϋg�󅹦�؀�v'Tv'��ن��a�@�$���q#S|üDx	R�z�Hp�ޅ`%�?q��_,�!����F|�*�����9F0Mw����u�u�w�Ƶ>��	l���D����}�e�n;�I�*������?IN59`R'(QE�����5J�<۪�^����DHJKF�v�[S}o�t`�#��|,7��k.S!�A�$�u����E�|E�Uȶo �b�26/u�
�[�P�tu��]} �3��;�	�}������+��q�eؼ����������9`K�H�99	BQ�a����rZ��E�FN�US'�)�t�s��GYHZ��j�@Ep8�m�n�{���C~�ӭ6�~C�v�I���T�
3)�4��s��%����[���^� i=lS�9��S�
���o�װ�@���X���Mf�Ʀ��O�����[w�N�v|�ڊj���#8�d�!k%$a}�6�;�i�,i�!C֭���X���� {�Ta��7˾�$?����W�R��AΕ���ef���H`06C��>�bn�"�<q�%�1�p�bDX�\�Ɏ��8���W�P��<�|�/�Z7���ą �����>��}��4��!����P������o��	F��Mw��uu��X,�88�5�i޾�cfIs�"-x@`07�T��Z�G�� �#���~�m_��T^b���Rg��_Cs��m�A�f(��继G�*Ქ��{�w~� k���M�̆ {D�KY��+�L����'9Ze%�#�ۯ������%֞��|�4IH�G�@��y~\⎛4����mp�r&vGƫ!,���"^r�
�f�դ����Y���(M(&Vo�ncL�Ғ�~i}�Т�*�ۃ�J3rW�P�+���\�����|v)pU�r�"��s����7m�w�H��y�<�Nvn.���*�;���y5W+�e�x:4KH胝�p��8.b�����jJ�s1�JNn�	��~r#x���_��Ax	�o��[�$���b�nDM֢��9�%��3[AU6l|�B�{�}T��Tx)�N�*�@\s��U`~���a �����I׈�h���c�0�YS��o~������?��|J�����^�n��T@��ϪO�
4���g���|�~ڢ��q���@^]�!�P���`+R:e�K!�?�5���E��xuQ� ��*�!��] (pi�t,�֤�4& ��zk��]Bw�R2���X�c��jlbo�ѿ˿�r����SDt�il��Y�t�N+��59e0�1^;��}>\J#O���p�a�Uk����CV�G��ҊP�:K/��e����P+�*ׄ������ֲ^�aֺ�7�6�GŌab�0Ъ�̽�>��2�	����z�+\'.���Ź,A���IaR�G(X|�2(��٫�������7�r�K��6�-��갲m}�c�g��oħ��A�Z��ՂD��^��j�`#ζ F~�_��b�@��k�	���~Nש���Pi��8�+��ey����@�.��0V޵�oJĥ����� 2�c���	4�E�����Qq�SdQHOF����r����T!��9ed�`��4��,�BS9X(�۲�Ŧ�^��Mr�8��{.�\3�š�M��=Q�[����ZCZ.|r�-�=�3a�+�
$���$�g���B��Z�x�@��y����<k͙/|ỿ�����W>��"/�u:W=K@��Hm�8��e��x�U�-lL�LL�KU�0�I�,Ts ʛ���)�����_�X��=n���`E������s����������s7��K �Lov�����J���e�M,�{�in���}?*�/]=�T����������G�'_&�m������.Bg�,ъd�+�Rj.���}��M��.ּ����89�a��;ݩ�*N�ʝ+W[w�n�Y���� �M�h�tm� ��5A*6J��i�m�O���3R9kf��b?-��N��b�{E���N^l���U��>��*y�;�y:��j1��'zD�2̖�� S#�F+]�D���o�bw�֬��Y���K�F�ϙQZ��Ҫ�,�0╶K]��Ֆ��EK;��M)W�%�+��NG�i���Ҍj�����]�@�.�V)z�G��N����S6A��ז���B�@v��s����\�W���5t���|���Q܉�;u$�`��"۫�S��I`�+����愰]w��/�u�N$����]�C0�L������i�~�Etb����0�_��5đ�����6SS'ǩ[m;a���&�VO��]��(�啣5U�<�z��O�F �Z�;���5H����}��c&�(�7K�Dy�Q��A����|Y�?M�h�]��]�aT���.k@tQ7�Hս���!��hڙJ@��tMyj�~���� ���{^U�4`}F]M��Җ8q!a����]<h����.]�}]�q���G �ܑy��c��2���&Z����!�!;OB�M��rMR8��|@6/H1��&�ϐ��_���=x7f^�w�11������ܓ���8���ɯ�5���-�n\��R`"�a��6��X����xJ��A��J���J��e&G3�/ӆbё(q�Ͷ�_�8��i�S��Z�b�:Ӭ>�ޜ�B,_ﾶ�GIϗf�\W7��MV/]k�G}xh'����!�"U{�s�Gną!%�w�M�A"����B����\��#��Νl�R;��ouGSӦ�ŕ�İ*�GP�-���D#.�nD9N��}L�@�:����<|?���ӗ_�f��P���G~���K)�?צ�Jg����&��Y+�	�#b�7O�[��u��an/�
.H /�bx�U3�C���Ԑ�\�eC���ʉ ~mJyx���X��_��
(����s����p��l�蟇�s߇��c�C�KAx���-�x֓�#o��p(瘁Zr��>�B�F��r�������)�����0���<H��1� 7��� K0�Y?�iV�&�4�n��o`1�$îg���)����#5���?OX�xdd�&͗���w�Č���A�g욍��|I���ׄ��e7&�#���+~�$D�cު�W�C�]�5�۝ SZ���`�۱�"V����␙�F��(����ް��qbזW��vg��)*EFY�?!�:�Zq����\�V��1�|��B�E%���ڝOimq����?�w�]�UA�Zrm���@ċ���!�-��<���3ޡ�� w���'B]ggW���:�3��Q�Mz>1\9�GT*�P���+�S%}�d%R���^�N���8~
n���UO2�۲bo����;��C��{����O�YM斏�,�½�)H�b���\�X�mZv���q����o���M���t�ҚI����逘�炦w����&�\j}��`"ɍi�r1�>}B�� ��Sw{K�9>��sb�It��?J�Y�cvs���q�XJ�iS�:�^mЀ��>,����{�zH��Eo&�,Ɂ(y1������2|n�f`���1��������O�­v�,ب*�0�I5.�=	n0���8D1���)��.��V�\�ͱ�����U�B�N(����Ş�� �P�����}|�}�Aum܄��%j68��ً5�����1�v(�w��5�3A.P��'/\`��^A�s.e���A�V�zG������j�zt|�����H�]�c�F����ۥd�T�-�:��f�*Պ��ֱ>�yϕ_��ؓi��MQE٤I1by��'ZDk��y��i�%��k�0�C}�?�gA�{�����E9,�~v�<cV����ͭ�,��Iхvvw�"�c�����Xa���t�ڶ��7�[B�h�@�Ã��#�$����L�U��b�q������!���G�*�w�-���y���^���`�څ�����~2��u$���>�T	�ڧ{��>s�'|�b��
ǑMZ��d�R}�Ě�10z��y�>״������4z_��|![h�"�=��:�J����I����ڿ��6��X���Z��������]_�ɽ�g2�Vh�+ʑ�%���]P-���4�6��-8��Gd��s����M\�N��(koG���$���jCdM���V�ϡ\e�GG����_0��l.8�~����<�$H$4�V�N�b읬��&���ʹ,Ƕ)N�88/�������Z��ú7_����}���d?R���T��N�ԉ���b���'�>�w��ݔƒ� vV(߷90J����/�$l�(u������꧛����IO,��&�Ʉ�/�琿���\��(s�Q�RN�ء�y�����l8���o#���<���P�P��>Kު�N�lDy��ҵR?�h���n�
Bkpk��~��L���TT�{�ې�ג���{FT>���M�(�t-��#��sȪR�����x'.�.,*��|h�z����eܾq8K�+7�p?�h�`F��N*`��By����Den%Zh��,�
|�����V����Y=z����#*d�,/�����M2(�	�g�I"�M��C����%���wA4����d��#(�ѷ�m��/Ʋ���6��#�����Ru��Ø��e\/3�K%�����C��5v�a�{�f���qU�L�Q��LC�^����G1f�A�jʡ����qyLz9�`�:���oC���np�����[4��-�SmzPHW9���l�32s�.kԠ�2�n	�)W�u�cu��&s��k����1�l�P`ey܃"��ࣽ�wBM��`��Y6ʔ�7S�-�AhӘJP��r�5��G�\�	0�eAZ@β�>oo;��2JƔ p�]�I~���RQ$��'f׽�*7�\tT������i+W����%s�`� ﻍ�;Q:�]�]x��K���M��&W?5*T4o�N�4 ��\�Bp�z���] ��H�j�gMhg�B���W��M����,;x5�cU��okx���(giP�+*\qb)���P�49�qpn}꘹���
� ����)�(��xZe�%D��u���Fe�KF�ċ� �������O�%�BY���w����x��cP�Ń��A�Yim��h3H����|}7�Os杖�ݤc��ς��LylM�w���D�KE��h��b��/[8�t���<�`i�����Ci��jx���2�֯�Gy�^�J¸-�KB��U3����'��*�A=r�<j�s�Egכ*!�l�3h�6rZ�������3��K� ����Aש(&���:��y gT9�X���/
�	g�Wb�k�~-��y��=�7>��JYҤad�� D
!��',��f,Ɂ�Jm�rv\���a]O��;X�0����Ѻ�l�L��X�A���b���3US,<y[�=�������=gq����D���ej��Yo���Pҟ?�>O�"eD�MP������&�x!U�̂���S<���5���]�	��>`���KobP>����Ú��Q���RT���@���<��sSy/A�O�,��X�p?�a(��x\�9οv�W���sH}�i|���U��
�@Xx<�S�5��1oTo<m�A�Z�����T�X}�լ'ʝ���--��?��O&6�f����!�M>�"��Y�]/��j�q;�d�Zl�����[���[[���Q)�In����~7�%JJ��kr���yd��mȽV&���Th���}�������R��"������t+��t�r���ky)��F}#S��H�9�2�k�\�g.C'x��B9�ذ�L</٣(�q����>w'}	��;|d+A[�o1vdt�y�ߡ�i��a��By,�`AnfJ���;>5h�^�6���ŭ�7k�P�;���*���Pe.��8H��6I��xm�#��������CQ܀@6z(8�m�3i���s)��T%�W���ߦ,o;�&�9,�
��%���>?��
���$�@�y٬�r{Kß��i����U�����Շ�^��?/U 7�E�99�n���}��|	'�z�����dP|�PG�A�?їȊ�%�]h��tMv�{�<U����
T��g��U�)�C8��I�N�
 �6��e�s!��j#c�6h��h����C�C~*2f/+�D,�3����{p�ǃ�		�����������\39�?��ֽ���5lФ�p���ŧ�y�Mx����b�f-�=�[��v��PlH ����~�_�R�';k�R>'+��T�K�>'#l�6���!0�oBm�p�g?̕���Ĩ���Q�1�ʿߌ*�$�;���/8��Vb��~AN�RZ��6�DU����c���rS��i��rF���{ْev��Z�Cm�x�e�d�Jiy�- @־��c
߿�h�վ� t�g0�\ꩦ|�45�o^��1��l��I��qe@���ݛXN�j@E^"�v\��������ֿ ��7Q�[g���{Bi+_��R^�VҴX�B[h�!;(iZX��Y�Fz �+��JH���PNgK��*�F{�KI�.�oC�.�`)*�"�θb;�v���\��f-.����ޓ�ҡM��!���e��P�"neW�d� .��x�S���^�LB�ƛm`�L%{��rVf�.�s#e��y�]8��w������2��6�� ��{�$N;� ��?Շ��-�^��Y�py\�ɺƦo��d�]6���x\���(�ȟ6��^H�x:���Glk��������	�]?�&�*ja�D����p��RO�Z��v�&�u(�L%x��&��U
��ѣ��L2�|E��oweZ�����Q��i�i ��+�J
Wy�tH2���NW�er����V�ߟ����/x�V�g4j���˳c���;�`�	��}g���n���!cpʖ����+N"Y�q�p(R�nP������k���X���)��Π.���َ�̈��ܰ��NĚ~�4'�,P�(����03�����n^*=Q9����m����y�RXj�s����I����&*hO}�g �Gn̾ў�_��
��U'��c�Υؓ��Ը�eP�
��G�Oơ��^�ল1d��	@�ɻ���YY�e��jԊ)=�x�ڷ��xx�	^n9�恃U�'��w�	�F2�-�%܍x�=�I� ���Xl���V F[6�����b����yo������n;As��~�-��!�%y.QcV@�G3����Bӌ�񔦇>a)���y�9D;P@2F9�<C�#.2��q�c-N����w��h]��8�����`mNy��:��������Mى�g�I?�f���GS)��ON>��`1WN�('������d���ۂ�L�x��K�"���Z��3C]�g�:�GD��� KP8�ɻ�!�85���ʁ�\ t��e!ȥF����H}�}|侽H��*�`�����<æ�h���P�~�c��	��A������L�YY��g���*yk��^@���TV�l��%Iy+%�>�#��1w�_O([<��[��标P�\{��=3�,Y�#0MҔk�o�\��t�*�d�Fz,e7}3Zڥ��|g)pe�!�n�������垠2�U�sb��%��
���3�'�3d�/�pn�x�����"n:`kt��ʃD�Lpֵ�>�j�����Ã�&o�GS����݅��ӛ�7W�6�=m~�A�W�K矉.�51�-��yzB�-s��������"�������"#��4��ND�A'5�����O�uC:�� �X^�%١�����'TA���Pn����KOe��cN����{�6�#�bZZ���x�OvX��|�/���F�*����df1 �V��*�R�~���׹~���q�Q�{P���fȐ[���E�Y��$��ģ�̨���Q`�\����g�Q>/7���Ɛ�Y�2���
�@��$��kt'��S���	��6Zw�e]��bHBRD��~z��NHbe8�({�BPH}�^#����+s����yx^�l�U�L���^���%�+��b�a1� �����(���E�R�H�/�|�/��u�)���y=���_�t3/�'�Z~oCzȏ�O�|�i��#��7�H�F����.�&�_oOA(��vf�"�lַ(Qp��?�y��G��Q����%�oP"~%r���K�!=vÚ�����v}�@�y�޻|�����3TK9�dχ���F_�bT���b-0���=��I�zK٧�1V��u`�$J,d�q��Ժ[Yf���5,Yy��-���L�`C��^3�ڍ
<D�۠���,v������t�|�Ir�#��!�X����7�bF^R�@�����#G]ï�2��̯�lsQZ{�'a����7��M�G'�cR�:	��Sߪh�׎�*n:D�~�+֭�N��>��NL�ƀW�8�����bl���_�>�8R���=��v�s�i*z�P�I�0!��I�l^nU��%��/@�fFa��M-MWK�Q7 Ӱ�S��3L�'֨� ���f��kD��i�͆��1�b�D�Ƿ���bǔ�
�_v���DZ�?�G�|g����ݏ5h�OL^�l�?�Ht<��x�8�d�����>��/_k!�
GH��{�9�������Y�VP.�/[���3��Zu@�rƎ l�v|P�`S{I��b�8di��g��'m��j�.f��}Q���F7�~uD �V�`��4�x%�7r�:�)�#�C�F�����fW֧$Sp�,�!8�7�(BqK���^���^/Pכ{vI�p����x�X
|}^�K�7|Y�׫�A|W|�P�Y�t=�L���ʗ��<�fe�+찳�p _�/rlr%�{���������6Kl��ޣ��8�8i�c����I��c��g�3��|�]Hŉ���i�i#&�)x�Z��
aݸ�z��ґ�4�4�n���z3���K#+���=[xf�<�"n(Oqs�k��M��� ->�U�f�~;��y�%h }'_��p�T9�2���c��$����x�&޵0Ļ�g�FJ=��L�|�x%v�����	��_B�'3�����qd�ЫU��'�	��>#�)�̛4͎�%K^�Uff���6O�^Ȍbll��Vs��CUF�X�s�i0��1��W*Qf|ڟ��A`ˋ7WLa�����r��kq� ����\��͊"�3$DS�ޚ�7��+�$0��)Ox�g�Q�AJ�SG�=��{�U��������o�Y���}Ė'�֋\<E��6����n��-?n���5i_D�˒G���E�P�&��&M�/��Fs��{kS�ʖG	 ̾ߎh��G�ZR���-���/���ٮ�f�:� ��=$}E�$:7��T�i%fJ
�/t�'���	ZY�������po�+/��_�r���=�a3<�
1њD������g�v�7��>(�0!/�_���)�-�B5���:&D����#O��am�nE!Ȣv��w��O�]m��S����Yk�M�'t�E\�<H2�`ȕx?9�@!Ӭ9�PP��n���v�y8 ��_rVZ)�!��Wd)�?x�nOH�Xͫ=">]ʊ��\�s�Pv���p/.��j�3�(\���6w��]��/2�%����>	��d�8��R��5>�����6n�C�#%P����o�9Q���C�~~姧�u�]�sN�"�o0!^ł���ӁSfeߚ��a�3�sn�a�9g�2�[�VX*��Ar°�V ���*A��] �J�fOH��ߛR�2\
um��},���8ǎ$_�l�y�=)[�dN8!��<@��@t� Y�5)���x����q�޽�5K\M2ȧg*�H�&s�v��_s�����P��FX�#�[U�m:�@%!���HVOiDޭ�S��<�e������u�s����x�?/�PI�xl��� ��T3�=w���7Bm�v:�����K,�ryW �S��v& z��%fY��rU�i͌���&8Y��۶@Ia��!][�,�5����$��z��I���K�'�-�3l���:BCN�"�O�6=�m����ό#�����{�E~���L �ĜV�X��u�uK�Ce���� V�|���J�)�/����U�����m�x[�}�ok�=W>�L[*�����k��4�4������|M!vC"3���_GWW��Sރ�<P�q����-g.L~��*a�jB�}�Gc*�����_����0��:���2Y*i��u�~<=�^°��C_���Ղ�Z"΂
|�������˹@��>1��A�2ű�YI�[j�eJ����Y"�~��!��� Q��=x[������D��D�\Hݔ�6�#�R"��c�����R�瞧	_�l����J�� ���%;{M�ه�+FeQ��(�b��Eňu��V� �M��4�8P��:՝$r���c ������C��o��8_�X�(�Z�������LC���@����!�u�.t��Q�߄��F9Pb�)��{�|��Ui����v�V��&��3ٙyk皿�,�T�+P��f��h��尯`�
߳�/9��Y��T�QQi:t��t�R����J�D�FP@z���4���.$R�I���K )�%|�������9���^k����$���ah>%~�`z�81�Zky�mCb�S�A"�&��Q�}��X�s�B���c:da6�;'���	仁r&_�mtZ i��y�R��tz�oyNocNCE �����N�����qˮ�.Q�2K��f���wXL�$�/���(	����fs�ly����nN���f��~��wVw�3V�_T��$Fj(㽰�F�}m�/era�؉�e�iٝy.�ͽ�]ߜ�nU��Tjr*�;�poS{�ݑ�,�w��o��L��>���������}󻚝�E=~���ۣ Z�Ƴ�?�[�	� {Չ����P�v��w�l�e?�Z�B��/dKҺ�����q�3%G>�6Ȓ��-z�7��˔����������tlv��M���I<m[R��=����o�k��K�O����'L�z9+dO��o8H�.�3ջ�z��=9�� �읭�C)���d�5l�Md��UC��h`I���?�}��Pt���z��R�#�:'�1HU�[�����"�zI�xZ��K0�	�:�zݔ$]N���A�?��kj���=�K3DP�9kgae�'�<��#�t�}��6�@^�\ǵة\4�?Z����M�G40��mLU�koP�W�X�2���.m��ՅJ�o���U��	� �1"y��׋���?�j}�!�K�\^���BZ�4���� ��Y�>F�m<���u]��<ژ_G�����;x٫//
�uxt�4�M�7}����0�Y!@�yc�Vrd�~i������_��kpEs(̭r~~K��Y�sW_�����{���f^xBK�(�e�[r-��� VP�fbt��ѩO�]���
'
K���Ej�k��#}�>$f� ��F E\��lz���6��|�Ҋ���������l/U�\�NC{{��a�5ϛ<����n|%������$���"_�|UsW@���[�z��>��X©P���`��M��ȫ� :�#��'��o^�	�Ni���at]քpw �/!�L�z4}��oQ�O�C��e�5Wia����A��n�Pś7 �� 󰽠gD��b{�A+X�k̎�*���N
��C��=!��˦�b~�$������5���߆���9Z���ё m�ٌ�[X
�������gՏ�`��<�M	�:DA�-�N�7q.�� Ct�\[�����!�z��m*v�T<|N{��7=֓�ڔ�Jo*����!x����E��[��~F�d�t=RV(;�!���:���D7���j�<*	���Y؞A{d�8�R�~�pu����hQg$�iP�椞
		�X�G��
��L�b0y��-��fZ�]�c��7�e�e���ʓ���̲ԯ�K�z�)��R�%oٖٴ��#?�U,���o>���.�Q�W�K��������@Q�5�X-�\�ǲƵ40�]�R�s��,��4A��IC�� ���~G�������4Z�}���PM�:#p8�R���gb���F��?��oԤ-
���M�O���Z�X4��I�g:+��ku���V��(��[�M���Wy&��y��I��_��~��:&����R��n��u������j������Y�/�m��>=�6;��������+}�����i�u�^W�A�����4��Ѣ3玮(pe?Z'�u�-Ę�E�o�&&��BzA\Q./7�>�Q��%����΢���i@f{������7N4#Z�Sϐ�;��;���O�����DJ�?D�-X;���u��3�U���E=^N��P�j��'�g(ex��s��P�����@���L�/v>J���[D.�� <�X��I��b��̔%uH�S4A��-�@�;{���L�8��}'���I�����a&��()��+��.#N�࣏!�4�a�/H��d��j�L�+�JIg�*4t�0_dg���
��˂��9 �
5Mf�+E����=J}g�	��0��)�X��o��7�9Eu�eF5>t�������w��f�c�Iz�.躙�)��r����P�C���^0�����a~���x��pÉ���A���<A�[��'}`x����V�:y��n0/��5O�(�(Y���2�I`\�)���Oc�O���-�����⫱��,�!�~-v�h����3���h�_�|7 ���������7�`����}��л,��P��et>�IyK�11	3�rd��$�h3Lr�`�R���у�i��/�M	|{3�˳�������{S��9bO�Ob3���������&,o���Q;�Xqgv��A-/��~.�����F+5��l�k⽬����9/����Q
8�D������K�w����ţY�ާ~h�ʲ�(]�t�#�j�M3�Gދ΅sz���nM4�C�(\��;R��U�C��J�µ�tI�@1���hv�id��@��/�����ε�?_����Ӝ�n��#:5�g�^j��`V����eJw�� q��9,�M�r��}�yg�Tz�D3����w���N���e���۝����O���xa��Pe���<O���zD=[�e�S8t�`a��W(���j�q�z�4��B�f�L�&��J�֨�M"O���������J���A��[�o���K d@[���>T>|�f�%Y]?Kp�ZX+�-3 i�d`�\/i�\��*I�,�B��lG��	�{5�6k�WM����Q�'�(N�omW�X���_��Ԃ��5(Ri5�#��'V�?Ӵ\t�L.F�`Lۋ'zObRG��m�� �O��b�aԷ�������E�������s2!�"��Q4d�i�;"�^n�Ô�[i ��5=��p������dyI>kH,hKC�rڨR?�[����A��_�$J����L�&��P�Z2�Q,-������x�?TRx"��<�PTFwƽ�����?���,ZoC۲j��<�4���Eut�C�Z��?)IU�/�y�]����������8��[hlbR�%�j^v�� �W�c�:�^wnѥK�1|�N�{����THNb/>�E���n���p��i��W���؉��)�K�'W�[��v�GB8Ll����|��$]�2UP�����1Ǐ3*�3�wF\e7VZY�i�\���I� /�؉��@6���Qh����b���b��/C�ge���Uװmt����<��_P��+��b�{����0w/���oBL�w����
���f�U]��f輯�����BY�t��t��9[�� f�i���q�A,��w�УB~Ě��S��ƚ���޻ /��C�l�8輸� =� ��Ј�!D\J��*���TskQѤ�#
��X��t��Q܉����F,k3�T�W�0�D*��;� ��R���Q^���lʌ�@���_�!D	ǰ]��(ƲFF�B�u���;@�e�����*�s"�)c�'j�'R�2�f"v����Q=�Xg������'�����i16(�:���`��2
ڷf��Y���m��D	�ӎqNk����~:���r�����̪� ��>Ua/����d<�Rc���H4Bv��0�	�:�����؇��h�w�6=�>ZP�o���ਫ���,��sD����wg�S�`�U���_�W���$/��nx_^]g�s>��M]��@���bI\gQ'��,X�An��!)e	���x�.)���IN�ҙ�����5_�h:�
��5�g�M��J-���\u�t��*O���T�M�&~�K5�$r��} �T�A����@�j���Z����}��zNt�>����e�z#	���Z9e9�Y�]���N}��ÓL����u�	P��8���q>�?����nq����N��m�/��m��KK��0��C������1:�0�*`�8�JI��c��d�R���GZ�J�� �/������}����[�GY'@��������]�?�q?Ò^��T	�e���;��B6�\���2c�a��$�osA���x �Vs��`�3d#����)J��
5Q��_�S�bKt��s-���Y�,c-���'	?�Y)�z*���;~O��U��.�=�>��-�0�o�U_6e+(o����������j���J 1�[;�C�6J��I��;�b/U��M��fn�y�)h�8�)��GsU�b(�I�z���wO0���#��>��0��:�1�d
�QVo���<��J��0�?td���J1g�J��3~�^�Pzp[r,a��o�H��0��|�xM��Q���'+�d�Dae��w��Éw֙��S\��3�Bb���t���=	� �e�R:����[��0X��,����&��:�4��_>�ϴ1��+~���������-{���\�^}��%������a�;[q�Mާ��f��**�a�?EQ:V��@�gvg 	�'" ��~(#���yE/9?�t�t4��sW��I��(OP��,�Șڵ��9�c����h���X&Jd��7hꮻ���;�w���7-�{7�NU5��?�h�;ƃ�C�ט)�"�?\��.��o���+9"��x3�-p�e�P[+2w����Xǥ�EE�I�þ�Y��ׅ~j��3|m^C%/�������r}b{��鍛-�X�������@B�}��)U��j����
��~r�9;=s�L�Q
��}�P��p4�&��/6>y��
p����vX�"YD�Z�=�'P���WecT�.c�6g�zyE���\?ۺ�-jKVL��܋��W��:�w�H�?�w�u^"�xj�9e����+92O{t���sAa���+����gT�G)��~ "�t(��|~l�,���-D����W�v��M�Ã� ͋�u�e�k����	Ը�Gt���#m����[ya��6��K�!
AΜ�yNl5��R��E+-k���q�	��0��",F�o������3	$w���ZX?ؑ\�L.�v䎒��Q�;N��ʕ]�1[5kx.���~45�Z�-@8�r�/��o�u�A�����)\�e�٩.�d?�$��jO�!��v�;5
v�3��|�!����h�.KP@e�ak��Y0�3��y��dd/��=�|~�h"y����*�Y���5���ws���QY]TX��zC��m�[��V�tUO�8����fR�Dʹo9���O�	FH����`����[3�S�e�V���LQR�L �{����2i皩�cv�6C�'����{K�ۻ�u����U��l� ��U���,��{��XcO�~�!��!
!�D�H��խ�*P�Y{0�T+��K�zGO~����J�����n����K��&��o�bE@@/�
�a(�Ms JDw���%��z��M#��a�g��٫1C��+s�"{Zjy������O����
{C��${>�0�n��+]Yx��D���0�� C�Nkɦwd�Sr����:(DU�*����.O^���u�$ئ��Hs�A���&�b�_q��\��x9Y������?7����F��k�NlK�$`H�BRv��i���Iِ�t�~L|��o���Xߚ-�bj����r̱x.Q�R⚬�辡Ŧ)QH%�cY-�W�n��c%A��]�)d��p��_��9��#�{���1�uB��j^9�+?��g�wiP�M��	f�C]!9�'>�9+����[��S4I���VJ��˖̳T
옓�E��0[��G�Zԉ%N��yib�gG]�ǈ�-�Z��E'tT}�(�P��p�s^;���R�&*{���ÖV�y�����V�Iנr�FF��8��-d�:n��K�� ��^����>��ত-��9���7&16>y� ¯��P�5]x���ٵ �}�k����vRH��͜}�9P�/G��	�l�:<T=Φ���ߜ�h�������R�Q���3PR�E��kU�#��/��:���@6�c=�RO�q76�K�$_�U�"�U���L:(�6,�'	��s�[K)���JOJ�a4('K�E�b��2������
�£� ���lcR߉w�HH:�T�^�4�)�|}T{\��>\�ys�l��5�qF�SpW�%�f�['Q'3����$ϲ����'ӷQkQ\�6< xْɁRw*�A8���\;p�zy�D 053)�e��2����h
Y����B�G�?���Pa)��zP�Č�_t��N��ݚ�PlJ��*��p^�P���c�'� .����Ue�3�Q�k��2�I��V�5ڥ^v6w�z�r��;��v©������Gɑ>_��������M�)�j�o�����ܚ+���O)|��}����5I��(�xb)�@B ��L�p��,��r��.V^��0���+�am�݉x*������{n�F�߲��)E�\B���Ⱥ�>=��+ɛ�I�t F!���,�����8^a����̖�iϠ+\Ps�I�l���%6zA�45�N��2��#������-5J@SuH'�Y��B�vy�Z�+!
��@���oe�[�e���)�����h[�D�Џ��,���)�'�	{�'4g��]�1�i�ΙSAE��	~�x����DV����U���`�PjU�y���P?�� <��5о�9��?�؝��95��Ѳ#K9��-�&�����\�y�β�=~>��~��4�7�(-ǩ�q�9�f��[��^�e=����b�,<�����1Q�U�3�����̓i��(52��/f�_k��?cf&��y�Ƨu@��I��l0��oJ �������i�Xf�E֡+��V^�ᤗ+*���)m�@Ŗqmƪ����v�7ր$�B�S�}\l�RА
�ͽ�~8h��w�v�bo�m�w��n=���
�{���?�7�j��qG&Z��s-�S_�1���ǽ_��Dz�E�EA�V7+<H[��9v�l��
�f ըV��i�s:_�e���N�<��w�X�ǽ��j���A�֜.t���OposS*ң�y~��;���e��sV�6�țՆ�=�O�	�fB��l�d�����{K��C����� ���gƺ3���2]cV��Y�N8�D���>���W�n����)[��2�.A]��#)v�����
��/��=0lE�3})Hi�GDPLh/@�|�x�.���I��IFgA�X�����`�SE�=�U�Fy�qؙF�u;��}��}�L����P��PV�H�)�}=J���_���*��4Kɋ�B��^�+{Y^R/��[E��Z��Fl������d�,�'�w����2���ki��,P��w��6*$��#�i$*q)"���z�?[X���&�S2�%~�{غ��KI61�n�6wV��������.�����V[7ބ�f��E�	@�қ��!��Lg�?!uPG���di�q��o�AS@;3�Hac/g:$z��r�ϻ�����$~X������(�n���V�gp�H�(��3�
j��
��AG��ӄ}�XpEG�L�E���=��&��T<�iX�!��	EA����.d-l�^e�z6H�.
�[���o��U��2�/���@���F�n�>����4��K��8f�2�s�=�VY����i�KA�C ��ӥ��7��Q3aSR�c���
0&O4V�q�� D߄ڜ�����*��������ד ���Е�:5�����2��j�BP��KΣ����;[oR���'�uzԦ�͚��(u2fG���q	�EX<��{Z��� �j�e�G�.% ��Iv����;ң"XH����h[�e֝1�tk�S�p�::�ߪ?�X[�)od��_߅&Ph����6�m�#�[!����Xhp]n��^�%V���Gx�ᶽ�_-���.p%6�ڢ����p���i�S�V���[:�	\s駷X=�)�J?jQ�5�� ��\��1��
��#\�b��qɠ��Y���d0-���X�߂~�5a����̭��M��1���NvQ��ٿ~�9 �ײ�;,�%�i-��
j�u�bs2��ٶ�v�O���d��O(���?��kl{3U5�p5�]0����T��|Cgr�=��{�JƦ��{:r��˪��ݹ�i�)h�}́x��EY��0���zǎ�L��%Yc���_[]��p��%<��0%:�+��V]��/}�!�G5Z��i��N�x�`�9�#w��Y�d�	�'6���7p,����;���jɴ�T�v�y5	��̪�	�qăE���h �����]��� i����=_Y��"��T>�%?�v�Wm3��c�fb 񯓎�����������0�d`m�f��k�������H$'��Gc�g�u��Y��iOj��ɻ�#}Z4�%�>o��M�R��71õ#�A����-@d����	���-���&��t:'����2�[�I?��grd��o=��H���Z��ђ���h��K����E�0�7�$+�4��E�-V ���~:.W�2x���	u�������u�%4�
���)M�ΥQ�'lv�)s��ƻ%d�l�hsL��=&:m=��������}�&�->bxL�bטC�jNH�kvώ���+�_+)����c�QZ�=N� 9�!�8M������������v�#\�%+o�����8k�ԩIq�R��A��A<1�=�9�b�*k&����G^�N����������fV:��{L����@F������'z��­p`J���9_�N�]w}m��|��7[~Wa��W5��2&��GU��|�/{q�Y3_* �g�`��'��>Q��nVv[���t(O�%:�i:1�S�߮��N�	�����8�
��X򧝯1$��\�5��lk�����}���_���q@�ݦ���A�oQ����� �2=��S`v0]��;�3L0��6�x �A�R�Y`�d��3>�A�|��7��3��%��1h��:��kwxBk�ѿ��Z��+x�3������lp�Nd���24#�x�]�Ɇ�6Y��D�T�pl�E�{��d�Z'b���������;z��T\��ʻ�'��?� 0a^�eA���Uh�O��4�3����`k��{�9�Ԗ�q_jF�� �2'�
�%�'�Td��jE�|F駟wm8��7��~R���ʞ�㑺r���Ɔ-�����~���|���M�-M'Kk�M�0��ޘ���z�WN���HW�瓝�K}gn��<�k���~�.������u��O�����XoZ�'�^@cG�J4A��!���-��j��N��A?oɣ�ki(�32��9_�y��O"M$�*	����񯙓&�Y}���qKͫ��2����pz��+%,7�����$hv�׹���e�A�%�;�*���!D�z�y�
LX������k���l>/.7苅���=MQ5���E�U���_����+��^tԜ�L�G��K��uy:7�?(ނuE�D)��5f�v�ǉ}��J���t���5�ܑp���[�vhe���M5wr�Xo�O�����'�9���'J��d���Z�j���ߑ_��s����̍wP�)p�V��.E`����'o�'d�����Չ��O��+M�_��v�	z�Aw!�g�ȋC&4�v�Ž���U�tq�sЗa�� MM������ms��<5M�c^O��=�ePg�ԝM�֟�3�T%���ى>�gA;r����_��oX��}Ŧ$��γK��xC	;B�h��9(�������}�/a,	g�)��(�(BW=w��ظA�D'9�ĜOwN�۪?Z���tG���L�h���갲��C7��[���Z���+*�%ɳ��+{U?�UW5�M5Oa�/�`//*�X�+z#��!8K�έ�1�j.{%.ٖ�x��܃l��F��z���#H��Q�~�56��.L����jD����l�Bu[�<�~��
���!D�T��\�g�tl͏�>^^2��2��Cᅁ�Y�r��@�Upߵ5�ݏM�l���(���c|ݧP}�
ԶG�@�X��M���W�waH�Eɷ��Ϊ�x��"]�N�~�i��	J�|�@.��N�"�=�mM0�nk^�����^�^<\ �a��O�_�Y"�����?� @q��ٽ��Y��**�9��b&��z*��nL�t`�@�{8�沝�?/����?��8�I�J<�1�A�\��
�J��6�k5�`*�t#��6���|n}}��I�5�����|�7����>��$��&(Qu�a��uh+h��=I�Ϙޠ�!�|
�oR.�B-�Q�C:-�C5 �r��WJ��=�d�*(����u%�Έ[7�շ�r�7P�0G���f\j��q��+�����keI���=u$]t@�h��
�X��b�����ݘ�ɝ>��g2���k����|3H�ZrE��1��c��߆WK����h���H���c"䌧�q!�)η��t�'��P^l�Z���R.ն�>O�F:��??����AKy�M�6��B��^��?-��n�$*:��L ؐ�yd����vA��#��,��i�D��f)�{Sv �k^a{�T6��V!�VGp��b���]\Й,?'p���=l��w{[�.c�Z��1��^K��"�tt/tQYWʍΦ�I��M�p�/H���!&�m�lg�'�"	����+� �:���F\���c[n����n[>�Q�\:u�5c�
��M~�N_h����|�?�F���an�\���N��ә�@P2?R�m�tx
&ٿ<��Bk)4�IOs��r@����:Jr!���Sk����$����������v�h����l�r�n�I�u�S��V��).��L��^��y�y���먨�*�Ç��$��~?Q�6�L�o+��A��H&�5�t����k�`'�u\D:h�u�l �z�� %J4J�u�����-pI��j֮��Ti��[���p�2�4�~D~�&b���Q �^?�:|�4:^����pL��Vq�ej�� !���03���z�������A#]��^'�\�.J ����|0�ͤJ�p����'{|`�7�H^=�4&�?.�p=�P��m{��t�-u���$�/{�{��j	�O��6�+b&L�S��Z�92�,2��Y-�b ��p'�����}FX�9��'?��qF�(�c_)�`�:y�#�^�A�8^�;y��
T�F�UX�]�@ �n��cVҗP��)u��4��:B���0y7��H��~�l{��U'ׁ��!�p(�{��UNI�i�ڟ���T��y2M�#�(D^���/�z��柘9�&b���Cמ���jo�$&��mN����)�Z˃J��������Zd����]"�A�q���fW��:s1	lÒhe��	�[�i�ʖn� b��:��F���XxV�F�*��3��g]^��rX�l�MdQ�����voU��w\�����Bo]��sVU6t����� �)/R
㩨@�0�dd �Y��e�f"�4���{Y0�h(f����m�]��ԥ�Bm��B�V��$�G�#��&��9���2�0ݸ�Ǣ�f ��׹�W��ֿ���G�L�%�]��d��G���7�����T :*�b�q}�.tfV�R�%鑝;%q �vzKw�۰=r�W��@�d1�U�n�!�V8\�K��P�S�����y�z�#{\�0���8پ!��]�&r�ӓ�0�1����B��
s���E�#�\�LU�dʲ��vܱf�:-uHBA�O��Ti�5��`�G1����}R�.\2�Sn��j�Bz�U�m9��_���A�n��B�#���p���������*y���"2��8�AF�Ic����_=;}�{fe����*'k���$odU!,!96���~x�o�T�����J؏-���~1��q:��5lվW"5���I�������%˝�5֕&���]|)��%�c�-%ک��I�X�纶��$�:�f�t��($:�v-
�N�d3�^�9h݋3�W+\�ؽ9��<��s���7^3,�]�ai*S'#1�	�����;�.�h���c(&��c��� ���ّ�Ed�!q�o#9g^�}��>p4HI�0�C�l�gK]����������o�Ő8c��S�l�In�=�[�gh��k�(�iV ���?8��@�Κ��{vƏ�o�.�|�����	��	Ҫ:�����j�2��x�[Ԣl�����j1[���W�����X��k8��mޥ�^:��EhQ��/D45`.�$+���d�L{�a��|va���yU��`=��x��$����2�z� � �	�Y��%�#��6�ug�j�ͦ$���`�b���g�3f��\qQU��V7�Y{>�5�oHU�]� o��e�h�����5�h�z҇���s��_��9<�c��9� ��H��[Ma*%�Sccr�GH�^EԿ���=��s��>���M�w�� �Ap�j���'�����ޫ�ݸ4�,�	�N�T(����%���c��k��t ���M�U˷:���49˖�ǡd5��@��)�J;���?�J ݗ��'y��B��u��]��r���-���p fQ�UȦ���A+�Z�jXi�I;� 8�]Tn�Wt�J1�1���b��^�g�D�7��[,�S����!59��$���"��}ش�Ŷe0���\n"�H�|���XzS}�^���$ɝ''?�II������8��R��,S������(kÝ�
+|�Vk�Z��!Q��T���,R���V@>1�ΐ~��[.t�Zx/�/Á���������D`�w�3���n_�w��x�p".�Ua���׃�lY�Å�n��-�����x�x�d"w4~Z������iT�˃o�uS@gu�#1N�{�ȁ��Cꄳ�C,NP̘�Cαrs
�D��j���4��j%��χA/Ӏ�-�@��Y��UB#�[�XG��f�����.A�yA	��웱����by�Dv�Ļ�*_���LsSs�WA�(��'�><����kY�pS�Ę�
>/��Gi�֢=���-�Ŝp �ZK�.#���LS��J�+Ie��g����� �a���5oyS»q�� rd��<	z��k��ˋ�}WҶ2&~@�W T��re�qG���%m�=��\�-9sd���.P� Օ����ݖ��˩���m��(`�A�7#���(���Ts�+����Ӡ����i'��%��_��\c�	�u��z?|pMb �{��|dgQ1��n�S�U�6�y�͡�KY���v�N>G"���W�^�0;!��[K^�]KlT*�$Q�z�O�Fl�5<)\1P�s(.�w���[8�Z���t�e���R���Ԯ�`w'#�,q����g��t��V?�4-�f��kr��NOP	��Vk�NP���(S"��pP�t%)L��Ȋ�&��d�'��}��7g+�Z�r���6��.B<t�ZS�\8k�9C�#�`G;���e��S��*�̇ug�d���TS�h�BL�Y0�'�3����KE�P7=XJe/��O��)���c���`����J��83�j�>��[9�M���]}�����﷒Fu�n�oap�Qԗ5A;��ih�Bm��{K��sU��<_�������X��V1
���Oj�7h�����plݛ:����Gm�n3'�ř�;�������k�j���y�g�`~d�*e����2UU��X�ޥ���(6��Nl�Ru�����c�鰙����,3�ga#��+�;��y�z���,0#�;O���ظe�L�Pp��[�v천ZX��lZ1`�@����;�!z��6\�6/J�c�@}+D隷�S3\�ރ�*��m�5��:J7�a��f�*��Y��۱�O\�:��绂�F��v��Ƶ�з��=`�#��|j��}i�l�ٰ��������r�����o �%|�� aw���f�&��ޠ�6�hԧ³<Et3{�䩅cej]tw�}��ݗ6�߁�O���	l����G�H��) �yx�:ha6�q���p�/Џx�ti����%�+C�㯝�RҰL��<��ԑݣ����3Ml:���*���ö(^��.(������_A���)x�����j��F��;����s��?���zg��R�0��d/δ�K��ޏ�� ��$�`i���=@}4��wBӔ��;�3]��uڥ�{a��>���(��`źϘ~��44��`�l L��-�$ @4�G^m0�	�?{pf�eZo��W0��:Tc�)3��RI�V�t���ã���.�:O��$P(��l��p%&{P	�$�X�h��O�h�����:,}=��\($Sf����4���ͱg�Mu���Y�Z�
�B\_���a�R�T�����C�>[���;S�.Â{M�����@ն�D`�#@!6&���^�ٟq��E��L|g��u�������G�m�#w긁����t~7>*��"�!�C�J�٠5�h�e"�d���u��nZ�P[���(Q��7�e�R"Oq9y��h)=.3��X�j���VaVCO,a��@�U��1����FW�~�fml����, y���\"����*/s�`@��?�����~���Ğ��E�l��5��i��y_�Z�[�[�Q{��i�`p�%�,��k��O�'�b�?�����m*�3���4�P��px�-cB�`�C%Y7��P.�6d���ii�d��Xa�j"f{.�2*�\�l!zl�@p�шPdȐ~��2U����d����+�r+\��J�7�'R�ɬ7# �ԅ���B� 3x�arwTF?�_u���3�5,��]���0��(_�V���l5&d�G>l"�#��~T�q���x���^5�x�n���m���Ym����rhu�r��h+�6�.��u���~ؿG%`=l���ƃ$VpE`X�r�6ݠ*N1K�h|�YV"[�U1���� ~5�~��G�T���;�;�o��Ȑi!$�Br�n��ka"�x,�u
��o�V����㋼A�!�bh�9�K���,����F-Dsv���@�?�a9�`a�[n�A�A+��������[�.K���$y`���T�RFD�8�a��:��瓅���'�ٰik\�y�ߴ���B���N�]�ĺӃ_�T��	��np���*^~�]�^hL���z�K��P�5��E_��8�!J#]�#%��Ŀ�Y
Ԕ�&A'�z~%��$���9�I5���zHt��Ϙ�b���)��%�G
]x���/|���Dfe�m�c��0x�jbx��<!��D�p�+z8h�$2��Cbh��@H� ɟ�޷�íd3"Τ�'��*z�:v�e��:����]��^�z��Bvu���(C��pF�*��d��*(s4��?;�	̅����Td����iNM��K��9��жTn	L��mY��
�L����)n�2��]y�T�׮S��(�h���#�m���[t0Iş�\��3XG<S���rRxI�^���.A��v�Md��]f�|�z%�3F��k(z�����q�D�-�nS�_e�]���D#�����-��o�{;����7,0����E���# ����!J�Wy�����
��'Bx�E�H>JC�d}�U݋��B\xۊ�SAPJ��FD�I�/�`r�5�.t�<��o��{�f���6	_빺H&�t�di,�L�V,���$�R���J�#r�P��Ece�6����LdW(:Ȁ<sj�:H�-�E�����������G��}'ipJ�WĻAS�k3Љ;��>�/���i9�;����~�_�e�7��T����e���Ag�Zz��C;�����U���Ȕ��|u�me|�r,���ɼ+��b�R���>��@PP䫣TM�X�>%� )p�&��[$�����bH��|���L� ���0��@940���t�e#���0���W�޴;�b�)n@C-�F�Zg�i����I��W� �ݘ�~�&��)1Zn0[D��L`��|�H��נD�� ��t�!W�l����*W%/ J+�~�������(�{j��z��}Q	p��ow �Z� '�33�`���FYafZb�[�)�5�ٺh��SB��"^�9%R��T��j�j'R:��l�D�c��(Q���������!4:�g����Z�� �2�\����:9�&��MGJ�&�j#��T��w%>�KW0�.��6|�h���?�O�P�&���֭]��~
���m���jP2Y�g �y�mn.��d=�`�]}
�S���5�_�#�ZX��΂U�֟cM�K���3u�'��{���֌fb��SnZ���[�=V ����d=,M���Æ1��pGȐ�)�x�e�4�њ��{�W�w�\�ϳ%��5���w7E���,2r*ѪE�m��l�d��rc�Ѱ��?��:n�I�z�����Lf��Y�ގ(�\�W�9��gU
��J&<�׮F�S�#Ug0�6�\3��YN�/�~u �"�d�`��SC�s�;����.�̺Ш��U��xS�h�\�H|^��^��޲�q��EYU�G����iN0Z�9��d����;
n���!��-�����Y;���ZN�b�˞������~F��+kpWB�m�o�`�� Q&m}�x����6�ݖ�h�^O�������}%�(�@�j��V�"t#ҟ(��f���0�(�r�dQ3�'��@䕧��U������|�y �-DΣ�te�E"'��K�%�/�af����z�ϛ~#$�!T9_�`�P8�i��r����)�XZ�8�8~H}�DR+l�yj�t=��˘�t�eg(]P����B��-��\��G���+̪���y��yǯգ�-lG	��Ô��U 	�B'��a��Ma1���'��'+LM~�3a�Kqw����%�3�����Ǒ
��ҧh`6'�`6��:?`
�Q%�������xXn
�� �����C
�&���n���JR̈́>dc��7��-eo-͏�n���5[���c�s�2��E�'C��ȏ��{2��EF�
�O٢��ږ���h�y��w�c�_��v���̢�5))��U�ɺ�6$����XM|�m_�L�/9�%�>�ɼeN�cr���w	o*úL�!d?��>�қ�z8���� t����W�@cQ�z��\_i�q�wj�.�[���t��8�>�BpdXsX���B�OV������sv�D>j��M)2*%#�:�Jb<��%@���ٲ�v��Ւ�v�у���/7���98����ߺ)XL�^;����� s�:ȧ���	�/!6-V�@�\v�z�ޕ��͂k��o˨� ��jD*b���vߙ6����P$�w�Q�A��ڻ��:KE,����hn�)YF+Y�]����ɴLG�6�N�չ���qth]Om�E�=������R��s9��1?b�)f�T�c��vy|�W3v�a7g���K�W��$�[�>ls��@�FCLE�#dlP�&_��27Z c��YH��8O������W���W;����f�v=���X��D����b|����u;Ѻi~�Z��R�n�ќ��V*,��g�꠲7)�3t6�����	��k�o�_-��~tR�h<�v�A�����'�	>�ڵ�}�g¥��~�~��X�<���ڙ�\�?.�r@a)Spٺ��#���\��񑢓��"B�NI����rt({ٳGQ����RYRɒE�=�n��,��>�샱o��{F������龯�u�^����|]�}߳��E�jVb@���'��=��q;���$=# ���̉�vLk��evy�h*`0�O8�g����6I�S�|���q�ļVK�6I�0���i��^a�ޭ����?NRʱ���	�����
��4.�0�7�&�k�:ה�T���z��қPC��tJ������x>��>�-���G��l�?����M#���.��"V����v+�۳���� O�+�x������1��ex��j��4a�Fe�������)G!�Ѷf	���:�v����!G�w̶p.S�K?M� �Q���"��@�_/��`�c"�\���ETje5�fs����?���KA�L��P�Dټ���/��q�t�餧�}~���E���~ �
Ц�� D��f�o�MI�/z<W�������Z�I��̲f�y�eT���lwΖ'eF��!�>�T���6w�N7����_�u����^�q+'�|�����`"\��:�9�������0KO����n�E���y7��u��v��S?iju�z��KL�^�y�z�v�Qc����l|cOu)��0�'��92:|����ޗ��S.QW�ٌ��L�.JT�Ga�/�[�A៩~�v�ZP�1宫>�[�3�,�H����ּǵ��1t���`Ƴ���
i��� ��c�Hy��{�� &�O46j@#�{!���9=̧<
�2}��9�>Lw�=j�R�Ҥ ��a�2�M]�G5�\>g&n�`��(p��.PO�o{9宽�c�Շ'A|��/���/#��E�f�$���β�?}.��n���l��)��GYK�-�G�dzKΣX���#R^��?4��j^a���u�b�ř���J�v�O>-���_�̒���j�L��S6��+r�:X"�!�5旑���Gj��wG.�t3\�����{5R���ܞK_�-B�&;Vg+�a�3U���hk�r�e�2�Y29aP���z�3���N�*�4��Ԟr� Z�$�q��c������%�6�s[��ɭ.�s�4�o�o�;�~�ϳuD.��Q(`K���+����.�%�Tunvx�T�'4�A�d�c��<��H���S�-{���j���e��<������^�}t?#c��n(�?m�G�QG��^��Cv~r;��Y�����N�E���I)�3��r�<υzS����A�_ab~����W�5h�t)�7�����~��2;�����%rȖiF")#֡��'�+[��Ҡm��j�ԙ6F����\z�_�F޲��-*��!EUBB�\��,e�^�wi7�ps1�O}���B�+4�?�a���Cآ�Y�X�_�2w �Q�3�Щqk�B����Ϛ���\y��&e�=�C>�m!���+�a櫕�zC����6�c��9>��`��u,ci0��ު�Sm�c���O�JwNk�	?``�7^Έ�\�;:��H*�k��ut�H!7�F7�ӕ��7�QS��V`�R��^�:��,���cH�g;��_�L޲M���;����`�y�f�߯m |��j�8� ���������c��Ģ�a�)<�'�N������ ��w�Gn�D���O?��U�Ö36��DM��B;b�,����=�m��td6�R-Â�3]ꮏ]Γ�y�W0��I�P�V�'��S�A �O(t�5�m�+w_��*�,��[1%�M��Ѝ�_Ɍ�@�8��c�(XϕGH�A�����8���@qN�w�c�i���%D�PU����
HJE_n%o�-����+��w�@�) [@GD�%�N��u.��R���.��µ��E��s1���Y�K��MN��`���3[N�W�(�S���w�H^wד݊��]j?��J�ln��K��(�Q�jU��m�ݕ�1���h���������X�09�ݗ�d�C(�=���[&%3lw0��l�"�����ur���7l����߹�c��|���(>��S�T�#ڮ�n�n[���n1�CrG�*f�j�8�.8���5���b}�8o�/���%��_݈R�6�L&��2ϼ'�R�2,�Xr��f�l�cҎ�S�%J5w/��Y�2;�[e�q���5-~H[T�㿟@�csP'�|����:|�͝�]x�A�k��CfԂ�3�W+Z�
��/��ܓp�M����om�=C)��(t�AD��O�<�U)#���lE6�p���/0��(X,��Ŗ���7��kn�q�z�� �`;E�+���;�������*�5mvc�
�!��&D�cu�r�/�SID��ݼ�Q�߷�׹>��U��F��'��?���$�z����[_����m��s~#�5ɋ�e3,�%��5��q�A���k5`p�� C/uq-S�oѨ�_G�e̯_�7�F�Z�/E�Ǣ:�~B`E�}R�I0�5�E��?�ڑ��Zj�wɻn�Av	��a��g���y��Su�f�^Bgz[@�Q�����2:I���i�k,�|0	/����1�8�����4��M�}�r�Y+�U�C����(�� �^5�������7�P��x6f|@�n�L��j�F��龃q�����+�-=J$�ti�:��Gh��k�$>'i�D��.�n�����ޖ���R(=��˭:��Y��6���Ȗb�!8ws�����#��`����Ʌ��͗7l*�gq^i���X]�b;�ǵ���2 N����+�3b��J:/�Y�8�`��0ܥj��hG}�(�ϋ��r��4�
D�� @Y�	�zˑM�ۉg�`����܄��ϴ��Νp�\e)

A(���Rs��xy�w�V}��x�6+de��LA�E]��b�V�<�׏��X$��fͫ�u�t=k�jϽa���7 �mnb���ڒ���wz�S$x���>giH���A�.�V\"t~C�\���e����'��%�2]q������SW*:��S6��U�5���-|H��or��_�.H�����
��E5Ϭ�����F��n.·^'d����zK��*��3��u�<�soAM˿=�g�: (�7��ߗ�/¹�X�-w�
#,A|#OEM����|�x�+�V�d��T�%���F����?Mi�Y��;�_��G�T����QVS+ܝRX$l�&���
�A��ԴV36�*x��G�_���_���TP7hud7����z橥��Xt�����Ոpa��-t�J4'k�26fo���V
��Tq�P| ��ss!|���`�+@��o:P��1W��9�� u�Ÿ��M+���-�}D��V"+@�	ـ��9`���o]2����߂�o��~6��K�X#�֬xJ��Aua�_�p��A<�Q(�@6���B�(��^�����Ÿ�e>c�>w0���?����K�Z��ѻ�v�K���<0��I%o�Yʮ:�$�vS?�L͍��0����ާ�7���$���t���t���S��Dg��գa��T�z��=]��K�����<,�ɬ<��ۏk'}�1�\n�J3���9�B��f������?<���Y�&h���H�Ǜ�b���Kݑ��֭�"�����١�.�����ذ��p�qWש���w̫�ӿ��7�����}t�RJ9�E�C�M�C�>^@����-`�)og9�`����W���g�@�n�pd�ޕXɱu��=�;��3�/s�ҹ4��Kqgh�����q0.��C�DK��~|K����G�7�_��8e1�Ov1���D�ׇ#�h�m��Z�5��GNF-dAo%�7��e��Dd�?�L�6����j0��ODy.��Z���
'�ۨ��1� Y��x�^P@�f��a�c�5n�H�_�$�m� ��,�Z���K=��Y�d�zc(I�k0N�������C��
c����B˩��W�˭�'�#����(�mV���T@��#���o�p;SQnc1���*v���W]�]���/s�����\Y�l�����������F��ㇳ� A���<M~�N�^�a�D�g�1S)t��e	�zJc�'��
W)[6ײ+=E�F�'D��vE+	������=M��������j���UR��;W�=�)�2�k4*�e�4ʂ��^D�VEF�f�?���1��9=\���h�ظ2j�Y]���J�\A��2.%��LL�\s(Y���}*ea���L-��=�_	�|�U�y�`x?Hu�./q��+���Z'+�I6Jo���!XB����i�Ն�����k�>M X�٣��4C��s� *>@��PWX��v3��Q2B*i����CD�bQ�� �p��RAi��(?2�x���K��U��#��4�m��ʁ�t��2����>	C^,�hh�b;'s�(@���������D9٠�N��.��z��=U���qVWB����h��҃b>����e����s�K/����洗��o=�v:��$v��wr&z�SJi6��\=��}�'�C��q������)|�����,���ۏGI�˻�}
���&��G�I#��,�����Dߖ��E#�o�#�#]1��y�2V��i�J�13xS.�A��g�Ұ��M��,�:���Ʉ�M�	���ȃ4�|؇AR�,O?�u�hkQ{� q�L����-�q�,׽�=/�jH �72��s1ȇ��dbV����f��T���ҹ�ֺW�@�e�4�;{޸t:�]s}634��p�ȫ����})��3 �"A�ܟ+_,�ה�>y�B�b���{��u��bj����~���&�(P�_����?�ʻL��8��kO���xZ���z����X����4�	>���​�&�1��NV�g�����2ͬv]��0r �&�%f���}`AR�,�r֧��>6��=,yW)U�fn�^$�*�zو��wB}|=�sAw�Y൏�8��Ct��8����ՠ�v�����\�w��﹗�>��l��#�_�����R%��1T�9���9y\���/���4�uKq�@����[�k�����Fs��}���|��JA��bV*5ũ(�5��;-��!;a��i�-~?���'B�1�\!o�s�69<�w���4�Z~׷��pާ�X�+�kx._wA�"Xk��I����5)~g@N<�+��kh=��1��)�e_j�2�y��K��A-����s�`�ݹ����	� @{� �� �{��$&��� ���5��:QLn5�G>�1Wo�yc�?E�c���p�hF��*\�����K�0r����R�y��v���R*���gy`����ē:��9�oB�#}�M&�щ;W&Ke��vJ0�.��6���P�7`�o�V���ɬ���R���2���~A{���T��"�>�J$&�ށl�g��@4)$&j��_"��h�!�A�kC}l��M@V����*�c*�U����*ZL�~*v��ZII8�`(k�����ޡ͑��AsP]������h���p���պQ.���-�Wqi�,�q]CWҒ OQ�^"_"�Dx�kw��,u�zD=���`����qX&�9����8�y���a�B��qB�:���U|��t���E��70@�e�(�9�S�a� �fG2U�l#��7>�9�����sEf�R˦�,�z�`��}� ��#�|��Ј�b��� �>eu9*��]Pv�wr��s����za��Z�z��P�WcYŌ���8�<p0c��N+:�LN�+v���g��g���Tmi�0^d�{3�Y��a�SL���I+�	�6,�]#��fI�'�o��d\��b8@/'GTV�&�6�'��0?!R8���Sf6��ٶ
�y�����[_��L���I=��Ȧ�B�'���(:Z�E~} �t�Y O�h֦z"C���̩_�����C/���X�+��!TCq�\640��z	�Qm���	+w�2\�޾}Sv�}4+�'�9O&R+7�W��7!P�+�r�'E��m�]%�ͻ 	I�k�v�\
.��B�F���	��E����aH���_\
�;�z��@,�������<n60]��~���p3'�/M2B&�_�=Ȟۨ-c��i40����w���=�FI�:���R)�\��{ݧn&�d�`�T�2|�}�O�>�*��߱�c-�O_������M� �:Y�����ά�8���tI�/���H�*��ĿM*eڞ�^E�_����cjFo��B����*��߾/Q�DJ� (�˺�l���^)�Lt�v�~�>��:E\��ƀ6z���x���b���`��T:��n	��U��2��A/�k!�5p�	\���m|������5jI�����B֕�]�ݟ5��$С@т��H�P���.e� H?d#��>�m{��}�K���ry��8�D�嫍OT�aG�$ř�+	��/�rB����gxh�6X�|�j���db�ξ��II��C�&Þh�� V�4-�j7V���7�����ů CB[;�F�%�Ȃ0ˊN�<���}�Ӵ�e}U�ؗ�6A�60[���}'�&��2��nN'A����#�e'�e����F���=�m��h���n���{�F�Zo����h�=��!�"�,��=�[��֤^޴)h�����E�1���3�k�*��[�m9T���}�g��ۀ޶h�w��7P���:/[���2���ֵ��X!��(��*��!�	BP���2޴~M�vxM�p#�8��W��^ؖ�����[����S�"т�qz$���j��O�?�-��3��̣�m�L�t��
],Xr�D�#*S�Tt ��!Y��lu�� f�~�²�Ke��+�>�,��"���Iqz�Ç��Y"�ȶԋ�=��j ���ҿ�������n�}�~Kp����߫l��M�+Y����d�kD�r�J�K�j�B.�HɯH9hD� ��7�����ؕ7�!QG����X3�h�Ek����so�/�8?�@�j�5�.�=�a�~.��2'ʹ�VIKM+�;�XX`��9Fj_�(�[�K�L7�(A�c���]��������q���Y�fr<��9" >���f[c9�������W��z(���)P^ +e���\����
0�F�ѵ�&~��0h8(?p�"Q���	ӸK>��2kv[�er�P]9P�E���bt�\n������8�L�9����˼G�4��� ��̓�^��w�Ӂ_���bS{���/�!T��Q@�({H_�m*0�}&�d�!\��2�o7�e�?����a3=�-q�$W�=��)�o+(�T�_n���htgV�I��4�p/�N��hdb���#��P�N�x�1�=������������Fs��bXz�����P_�n�K�_Sg�ꤵ��F�L�Y��t8�{�C�%��F���[��m���8uT'�̧D+=Z��'<ު*�Q�h����:�:x��f�oE�_7�3�F���m�����/��� �T��ܲ����Oc���<��%=0qU�64i�*�.��U��Z���OkRp��ı�c�֟ f��Oq���>L��J|ti��Hi%r@�BM%���q��#�S�e�\���(u�^ �n��>�{G�aVHd�ѻ��ب���Y���������4�=���Я-;������ʯ�M�A+Q��K���n�C���@��բ������J�Qf���I�9K���Ҳ�!.ݬ��ii���� ��.&̀��i�Q���2�%U\��_$m3�%.ޤ�H&��"(CnT�Y|"�}|�+��ÍGP'��S:���|l@�9��}��Oc�9�ٱH�:�g9U7�4�1\0j�.�����1��~����HL:]`��-��r�����h�C� dF��YK�n� �^#&�S~2#�H�@��S
"K�D�x7�FP���9o���혪�7�6?����nqP����@�z�|j��u��Ά$�$ ��˖� 2)#,��ihi�߃=������D�C#t�v�-m���;}UV������d�	*7}�V���@Gu���L�Ф�-Q`�3�PC�.¾�Z_����kU�7P���v�/�?����dYA�:	8����qF���	��`��*l{w+����Ä�ˍX$/�{�3��4Z�K�H���d�>̲%��_y2�TFJ����ͻ�nD�L\�y�%���ѭ�8����0����A�_� I�b�y���Q�Y�-Mu(��U�K�.���@�p�����L���SH���y�s�zg��?v�P!��1���+�PbCJ���B���1ɧ�s4�0�a�)w�w����Aփ�f�g��R������0�ˍ4D6_�+�l��x0�`��cNM���j�Yخ�a9;]���ϩ8j
̈�ݒ�uvD�>���[ίY\K�B�V�Ae-�g�8�A~R�H#���wV	H#��ns*�`�����/P��z25��vU%hUth�ߢ��5��K���@��h�����L�dl���~�F�>n|=�lA���n�""���~� ��٤�?�m�)b��~�r-�krI'��-F��r�z�E2��%[������cfv�֖A�~�kc7v+��-E�[���ܩW�ڶʉH//�-�O]�S��t���3�K"副^�ʣ	8�'�ћ����Y�Gp|�$��-ktڏ1�"���'�8@��aP~�*��p.���
� j�g"߁R%yjŬ�e�D�Q|�j�� AH��~��pA���Ud�2�y�ƕ䢲S�ܠ�W�q��U��}7�v�}�(�R-
/��uu�֠�ӏ�T.��&���uR񮸧5jLG/��<gY[�N��l�[�����p����B�ߍ'����t�t����nF���G��J"*�7�ɲw
�,����s�������ҵ.���2S���p�8�aL=X��^ʚ�*T��v3�u�nrlZz�����}��֊�E �4�3��&�7�6�a�'��hD���� %F��݂WWM+�L��:8	b��a��1�p��t��jL�u�8@����<��D�-����,��\!nCU\g�ˊ���n�����6?;z)G~k3�|R2N�����n�e�lnn��.	 �	����������bIx�zN�J)�l����	�y^�l�Ey]C��(<�׷8��"S|(R��T�c&�{?�eS[n���ԕ_,�E���A�Pޑ����.����(���:4bQܫ&�іp��ƪ�M���St,��e$�3�=��N2�J��[��&� x28K���y+h�roZJeg�{�� ?��+�t�}'�|�]��$���?��8�1���'8�ÿ�S�ڲ�������{����M)��e�m����T�	��i�W�"`���5/�ˎ�rzMGbvD���&��M1�B`�^
P�$̊� {��]�jr�������s魤�qs��Y�j$#Jp�{��~�.F��5�Ȇ�g�q}}/u��Y�3\ՇT��1{e;W�.�<8
)����w�V�P�:�n������G{b@/�1�� K�\.���7�Z�n����ś��8y:���IC^H���b���l��	�A��q���Go��d���=����W%���̬��ɑ���:"*�KY��/���I��.��A�����e��
-�(X&~4A��x�/ ��������I��E�5�IA=ݬu�c糼f�9�F�: �һl�Xv&�3���:�#���>�Jٳ����0���3b,��jg��N���̮e}g�HN:>p��C��Ⴣ]�?��Su�@�f8������̂�' |�^.ڂ~�ci%�����E��/��4��T��ڹ_}�͆���E��"�3J�\�
��&�����~�ř�X'���ZI�	��n���+~Bu����e�VdN���*'�+2.�9��(��󛻭�3��>ތgǦ���Xw�g ����k�F��8�ʤ��S'G�?��7����^���~klؖv�nǢo�I��La���ay�����8,��Rp�þtv�'<כ�B��7H�����D��A��Y{t���KX�2�t�a@���좠�3��� ��ۄ���~���� 3�K22t�䩿�֑������P�5�+��WR��N�*�(Q�O]{'��r�9&턵��i�I  a�J̨���/�O���ͷ)�5=��y:	���GV���G�`����é�WÇ�B6����P�V��4Aۚ^�V���:t�
�f!NO��y9ā��\�>8�̈�Χ
Ħ��DnE�׵1hm��T_򗗯;/�T�`Ķͭ24D>�Q�����S��%�k��
!J���.� ��&W�?�a�{��Sǎ꽠m�5|,��)/�} ����!!\_�i�����&�k�LE�C��Q4S���p(�������u=cg�*���5�@�j�u2��%8_&	'��E���U���������+x�H_�奢\��6f���=����Ow��R�[�`��L�L���������ja����X�0�Gٛ��t�}�����D@�_��~1c����4��w�p��R1�H6�P|9��ŷ9�:����
���2�1�)�vī�ߪ����^'����ö,�������ٻ�r���[sL��o��	��p�\���u��m�iz�<�KՇt`Y^�am�́�NhR$5����R����c�O���T��9Z���5Ȯ^�CqhI�Uh��ǌ&h)s��u|�ڠW���!%�U?'?b�a T��S59?�]�Z"*W�d�'�Z��JG��t����� ]� �t��ny"	��!h��`m�츇��x��N��境4k�,Y�EٺI��ub,;���?	�_�z�Bv��[:^��2K#�}!��X=lބ�����DKP���ڛd/�u����N��1MX�W".D�;A�|��z�z�>OM4��<�Is���,:S�m��e���M��^��Z�������p�4��?��o�2:g�@��QV���!�A���a*�H�EwYLJ*%J�%؅<2�ux�=�0�V����B�k�v-?x�L[��GW��uc8�V��IK?q�U�������>B`��r�o.�����7ސ�tI�[_҄Ž_�,���L%ORi�ut?b!�%xt�� �6��٭P����b喕�X[4:E����k$Mde�F���H�r�-���1M�da7�>#���vL �ی��z�gt����u�f��yc+���!��\[��"�
	�>iQ����H�Zx��LAZR+i� �1�o��S�Z����Az7��h�L�y*�D�}��R2X�$��j�߱�Dx�CN�5���障:��L(H�=���;:�`<3�QOc�,��ju��~d#g=b��E��(1���=���n_ �2�����=&ъ/{��
�v��%�ؓh�r�;���%�7˵��N4Z�H"��o����NB
m�M��` �]GЕ���wV�*�.uwll^5�yih�.���0X��\��9�l�~R�S�^��Kx;�!~$�ˠ⪇~%��9���d\	zT6���s;w,��
��E���#Q�|�f�T%$��v�Ukg�!�7�l����n��cs���g��9K+$�����Z���@F�����}c�����\_P5&o�g׃�מ.�O0�B%��l=�Y��Y�}��/Hݤ���6W������5��� ��5�}��wv"u����$1���J�Y��x��嬽,,�'�®~8��3E��j���{6�����xݻOH0�U����h�m�hjv���Jt��J��J����ĢB?-��q��A@��:i���3ke�ͽ��%���2Bq�pj�*2O9�QJ��@��!����f;@�֞��̮$���d7�Ӵ�\UZq��$����.�PP��_+,h0�SH��8Mq[TG"��l� ���}�nvW�5�������=�8���($���[�3��\4#�}e���Vf�f\�MR�{qx@�Hb6M��
kK��E���Bbg������h0�MŬ'W�N�'f l�C����y7�(�ÇW�)�5&��X��(�Y[�l� ��f��脲�L����Z~~\�}����m#���73ܼ�� �z6����.`����zC��;�4"��"�@�S�U�h����T���2�aJ3�hX�D|����bWh�I�;�V��-�J
���p�Y8K�ŏ��[��>h	"�{&(�͆JD I�6�[|��]��C6]I�h�[�y�"�J��������]b���o,=��d�ֻ�Nm1�u�n�9���mv��W�T��Ϸ��~�5_�7)���X��!ښ	@��a����J�N������u7L�v�s!Cy<E���QƮ!��֪�|�׬�/6�2Z�J�<�E�i��	�)��d ��i��^��LIj�>��AD7:�ۣ�o��M�p+G.��>����P	ShrЛ�J0�[j���ʢ]~���ZMa��A
�=���A3�E��F�S��yS3��*z5�K��������^�e��7:��N���:�J?L���f$m��a!�.z1����G��{�X��r�=�N�t���	~�ޓ9d��;:E�;������WJ�h������:0�����Z�]�`���Q��^�m��yr�1��&L9���.K�Бu73A`c��'�
�\�d��AE�>M@���2i^5tʜS���+t���w�R?2�&��2h�����N"na�xEd7�����bH"�'s��.2K*�2'��������[~+��׋ًk�#�\I=�����wj}b���azv���A)�Z���ď��}������Ȥ���U������Lkٳ�L���.}L���%�E�c{��}qI?�?>2���"�TG��Ql4/�0���ԅcz'hesMrQ�j�9G ~��-Ҷ��<ψ�xc"�7���-���LK+|����~У��Tg�� ��_�ȕ��ֶoR�n�OдŚhy)�h���i�%xd�L<cs����G7NsTf�r��	�r�H�7��(��h�unbHly3:��&��^g����F]R;eP�1�Ƅ�ݞ�@<�s�p�o�ȫ��*a�~/�������r����2U2�I � U�C=�*�X%�����p{,\�4
6淍w����k��a�6D���pU�( �������h��Jn�1u��}�"Q�����YAd��P �������{/�/�0���no���ޘ���6�2��9���ɧFV�����=]����~��cS��&EP�z�"a$@�{�E1(/%�N��6)�<8�e�k��=���Bï�}A��8��}0����ڪ��E����]��԰v�����9�PbE�ڵ����}�.jL:�ςu���Å_�=�q�@m�^���g�m`�-�qS�k��:�D v����`�T?G:;����sDn�(3�� 2(2i4{n���,�nL���^�^&%����O�a�1plE�֤�wޗ��	�g&-��t!U������_���"Qn4���O�U�!�,�-��T���s�ug&�en�vCR���I�0(�}A;��"/�#���{��%n�������!�Ud0������t�B@��f�����<�F��Y��%Gn����?ŀ�$畣aӄ�W���ȇ���������K3����}�ĸ���M����̍��\oB�cn�겾P�e���|���<͂8�	 ����UON��\h���$���(Y;������Ʀ^+ҫ�J������<�Q��Z��,5"�]�萼X"-�ދ|컼��f@Y|��H�i���<�x�wy�끑@�&t��q�-ټ�~6�[�O3���<V��	 �K۪�W�/��_�'�O�K��A�|�ė���qe�A����Q��"��"���=\v�q�a�FI�t��S��g�!(H�|C������+��d]����4-�9m5������Vq�s�Ʌ�1�l�?�{G��Bj0M(�hh{[���� �5W3Pӓ�Y~��"1��j\%��.=��1%��.� �ղN�5���2NK>BdxS�=&��A�(L�z,u��gb�n)!Y"4��S��<������
 ��IoZ�Ҍ;�Σ݆��r�m�ΔP����T��m'�����D|���lDj��R3���k�j2��$����ro�ĎS��pO�i������2?���\������L���Q8��vt��i-��i��e92j�;�0h{�攍����1
��L��O�p�pA�����J�}�^������ŉ��.��4\��y"j��Htw]����fr�_����Ї�N$M��ܦh�T��\�ۣ��nպ�q�'F�����d#9w��t^:�䇖�$y�mq�8S���z��eq�ɟ����@�م��+��dM�"��Չ$P���{Zh�#V����p����K�7 ;��FKq�u-����d@;&�Z��;W�$@]v�!\g�����Ҭ���E��l�vazMJ0ix�vl�U2����3�H�گGL������r��.u�z��֙d���,�` θxg��e׿����	|�ϧz�pĝ�-�GU�a� ���
萡3 3;�1�i.Rt�Vt��-���HM�'�*aT�!�^B�u��G#���?��ꮛn��j�'f�G?_����m$���$�k���6��"R��xzRg�*�L�s*�߫�Y:�O:�����:�:����`���N�	��~m����/�=�U"��J�"a9���\{�����\كA���
.{��s<�����/r�W���	�g�:�8X�Ӵn����N����Q'L���}*I���)��Դ�'6b���Lvxy��-B	Ǭ��16a6f��G��>,ɎL��BG��u�q�<J�s�A�R߁$��W�����s���Ҏ7�VH��`��D���,��+�^��M��p$vFTuo{�� ��h[��E�]�k�g�W��(�h�z,�V��~�>��p�K�z/0��*XV����1b��xR�[/�,�x��4��%��b��px�JL���Aڑ9HJ�k5�Rq���偓=�п?��%~Fڰk!֮�N� i�2o&��pm��v#L���Ո^�,t��\��R�#�_h�_��d�{�I�{�1���i� �r�qp��UU�q7�Hޫ�����T�_�NYH�Պ�9Ln�`�0�Z)�uz� �UTS��(�^�4§&���v@S�uI����[+ �����M���ݘ#�u���M� ��:��Qx3��st�7cy4�um�4
�-�$M�\�`m���Xl�vi�mnG��/ �Q$P����{�|$W�&����ߥ��8���Y�>���G�
�K�n h�
o�g�f�Q�Lw$�6m�=��ҏ�(?�m�]��q��g��~D��5��)���UN�������c�YX��|��*�w���CAXF��<s0eLڦ8���_�K���2c'ROF�<�� ��j��Ρ��`��)���ty,�ؙ�:�N����)���H��{� ��O`����FVr����\,���s��!a�|
���5�@'��T�{"�I���
�P��H���?���(�����c�Cɦ�Ȏ�Kd�ܖꢠ�-�A�F�<���Gpd{U�
i�?�H���9�&߳Ⱥ�PJb3,HB������v��d�V��}eiW(��!�)���6;�	Mo���$Ĕ E�=篆Y��[3:sg?�a�¯�̱�D��sJ܎��헋d�f��F���A�)�2ё&vg�|o��Sԩ�M$Z�Ў�N�X���I��X��.��3�)WO��b�^�"�4�U�� ��Z�t3�$w��@��&�,r)�l��{��b����A�{��n�A!`QQm${0�ݘ7�O���%��Â��*�5�C&�'/xP�z���-!�مI�G�����$yUpA.��4I_�Y�p��2��v��i�T��USZ���ad�P0���/�(R��_Z��Rm��d�5Q�I��o�љ��t��80�.]�w�� �d��1Dd��3�\s�IT!� �y�zBMG� ��/?L%��`7���hʧ�0u��GjS�����12Y6�äO�*���SW-&�w�&j;�����f�JB
ψ'Z_�a�~��y��κJ��VA� >�ON��_�^��:��� �1���k��1E.a6I7�}���d�M�]��k�J����Y��"��R@=$�9��l�^-���l�Õ�����dJ�a�(k�\����}m���:�$b�W��@itaG�S�(��&��r����CX�����qy����>'Sb�JGf1��|z��w7���%�G�^��	�s�p*q�A5h�=�H@np~ �i�l�x1��H���T�Y~��nPT�?�s�gb��'�`�������T�kU|h����@�R	2m c��r��4oJ6�D!�We]�W/]7��#�8���8ғ��_z-}�AY�mm����W@��^�k��Ouw�\������)�sq�����| xI�̿-�Ț!҆y�݀��.a�k�[tK=�����2���|2eE���jak_�*�ՎM�����~+nz���!R	����X���x�I*37wTUZm	���:F1���q�_���e���Ԥ^��|	"�un�a6	��ǀK�Q�K�M<��ї ��v�����e�{��G䮀S�d�������Wv��p�U�l��KMl5�v�赬Id�(z_��A'�� 
K߉������tKx�(\��	��.�(���P�yf%mᘯ���=�eP��&�v�h�ƠO�#oimOfu�j(W�k�_\8��醖 2+��Y�^�6���ď���OI<s�L���PɘYF�{_���o=%���E gG;u����8}�B��$8���H9��TL��?���w"Ի�N��s�B�Q��l&�qn�~�FL����&}�~�z��`w���p�U�R����5a*K�	��QL=���X�Y2
J�:f�����?�i!�k�a��.�O* �މ;��l�K%��+?� ߳�*��EE���
�M���"Jd��eZA���a�=��'�8W"��C̠�S�>;��tF�_�`��Dn�M�(Q�U���Iz`�u����`=�W4f�5��3����t4圖5@w��U�oq���i�D{@7{T�����ŮF9	z���Tʋ-P�&�f�@�p���>(�8i�^��O<� �	ϩ���4Pz5R�;�������iyz/r�4�x�n�Xd�Cq�T�V���1*��ƍ��6�1#������ts���`�(��qs<U�F�_�L�I
�����=/mz���~`�.7@�O$�M��0Z�h\��/$F�W?$�Dd�&w�uɟ%��f�qix�*��s�D�R��h���W߼�h�����K�
Zp�WGo����m��_,��k4�̘�0�f5���?��ʹҵ�rj�%�-��g��ۋ��'�N
�No�0S
�[�"��(5".� �h�|{<	z�wqs��^�	=tgmm�yiS+p\,���A`Ӵ���fg)���AV���Yd�Edc���,��O��ّ��=<�0��1:�T~��3�����(ĳ�3�0�'��������X��g�V�s)�gU��6��0�'�}Qd��e�}�x�Kv�;���G�jĻÓ�6��a���v��?�'E������$��`�uB#;�VFM�e��E��g\��,Q��$m��t}
�n%,5�a_��p���1K�
���Eo@�q�WA�1����B�tP'�x����`�Z)�gɝ��l�h���1'��V@p<uz�cT�]�|�������&�n���[�%�ֿ�RմPL��N� �'^�i�lf�����Np�ƎZ2�L���z�=VMŀ�9��4͂;S~����Y���!�͎�䃫�	yt1�"�B�T\�kW����q��+�|n�r��^��\��#�I|�l\�:.E?7X�*�F���Ƥd'е�[�ƽS��7��M}�y��H��S���<F�{]A�5ȑ'\�v�˩���a�*f=�j�N.� ��i���P��4��: �vU�%HfPl�R�5U�b���P�4oc��[ �g��a/����!���H�a+!�q	��O`8E�@��*�[���x��ਓ)X�4����+� j���N*s��b0������KN}�
��	(!V�;T0U���{�;���T�&����v��0���yW�[�ؕ��J��@$�d+�;��Ml�2��H ����]�qzl�ڍ����v�-O�QѨ���O7,sf�����;F�,�
~=mbi������Ș�fv�W!G�ߏE��뉓�uh|w�p�8��8��]�2��i�S!u������!Uә�g�
��#���PmH|�q xv"_L�Ɛ �i��]n�ٳ �H!�- �ȍ{M;po�ć�m��H%H�>��k�aw���t��0��?�ô��w,��z��Hg���&w&�w�쪠�X�"�!'%�:媨��gK��e%�8jV �#�,dy�@��%��m�{A�2��%��}�ڴ|@O�a�t���b~[��kzlUKa��M3{�Ew\�X�H��滛XG�O`B���F�p=��=h�J�y�<@|g�S��� ���d۹�b{\`]1�(�E��E]
7Vz�˱�`"��p�R�Xӛx���*�։G���7��j{��Ͻ��݊&��M�p�P���K!s)D�2�~)n*���B�(�tЕ$�☎1���}��{mq?߿�����Y{�z?���<{���J�q��
$��1��{�ا3��c���p٭0�-"��Ŝ<nd�*�
���n&��â���һ�q�J'I�D��[��r�+���<+�2���y�q�,��IK9�}v0;H�j�x/���ke���a<�@T�ǀ4t����H���Dl�ytA�F����i��K�_���n���
��v��<��<w�f�	�K-��c^�:3s�e>O�-J��@}���#僀�"Yݫ�W��i}#�,]�w#y���CO cU��l)�=/"����Z#�KRh��=nS#�Kg���Hg�n�����.JA�|ow`F��)��X�$a�%������Y��Lqe������a�T;�7���+����s��}�� LC���x��Tpj���)ɸ.L �Dc篽��b(�9JѶ�l�,J@�`���d�3vx��XW�0�����6�)��?�ꝱ�d�e�D�in�X^W�e��.p�z��Y>nzs ZM6�3��(8-Hϭ���-�˗�^��ܞ��$���Ci�zLa���Gk�����6ؔ�p��:m9*R_�ÿ]4G���$��mH͌۞����E�����Od�:�݄BI��*~r��[�B��Uc��?��!���ͷ�㸻^{"-�{��y��=7]��vM�l�������H�5��B�&�i�{��+}���'͆ߖ���X�Q^u���wv�䀯>Gm�l�.�������	�b��
�D'����:�3�[��`!����6�BU�n��b��B2 �!&I�I�T5�����М�?;~F�.}�ߥ�]��ťKr���-Ǜm����O�Q��t��7�����|�.Aݟ�X�<M:6�����j�3����F��+�+a&���5�d^=��~����~����~����~����_��px���2q�}z붡*�v��Nyz`�q/�R��'�TBJcz��nX.љ���e�BP���Mѧޭ����;]P_��Ks�nr5�r�T��!T�#��6U(\߾�\�;�r�o��S_Lԩ��_D�NX�>�~�#�F��1�+���W�e�.^��{}��tW��$�����i���E��7�s7R��M6���tä�Ͳ[��6{��:��ft�w��:)��me��O�ʋ3�Z�b٤�I�2���s	���!��]�	��L~�tdge�r4���}���|��ir��c���ϥi�!\�#������R�!{X�+KZ�-"��"|�O!Uo�NWN���+�5$�Vۧ��)�X������zݙP4�Ċ�՟���&z���I�����o�L
�N��6��1���뢻NyV��|�݌��\D�#i�����Â
�4��������7j�|#�`�(U�����TS�8��,+�	p����^��j��Mf:K�s�"*O��{�\�����,�lN.ڻ2�����17����U	3-��t�ͰuD��W!~q{T�b]�8}��t��8�Sy��y[p��;H��7�?ZڛHL}�{e�j:f:�a����c6`p!/ $�꤆lBf�\�b&՛�#I�.�N�h�+;얞a+$�۱�t7�������6�;�kxW��y*��
m��Vb�:_N�KԌ%���Va� ;�輀�y$YՖv��5���~9��q������&�g�>K�DJ����\y��F�<ƃ�w �|�r�����y��b)3<?G�� �H��K���y�Պ��Z��'@_�]����KcKB_a���-��Ѷ6»�]��0e���I_��d�l��q�lr>q��Y0��4�b@�f�m�Y������w0�.���f�,(��A5�z��jK�Js�؇2M|�m��H��Y�p�N&Q�������Dn�����[��z<��h���URr��J#�ave��6��u���S��V"�s9WR�隆�,���w)�J��nA�_�N�����͎��/���L��_1`�P�o�z�$x�JZ���#;_*����)�M^[��ۄQ��=��ApO���쭔�K9Cv�~#����=�1�BhJ�w��P��>�F�cv��)�Q�fD,�[�ˣw2賾=��8!�G�5q)k�J�d���:
���K3uw���gjD&�Y*��}��G����U.����ml�0nM���\$��_~Mz�M�o�z_�w-Z��Z�Wp�y��>�9����vY]�����W��sS�N�o2_P
�_*�]g� d��s��(���&,�qn~��a/��kZ'�J�{�N43	����l��n�o���'���φ�f!̓�m 7�X�±��ey���p8���Q��?��<({&T$���� �h�ؔx��b�d6F+�f����v��S�[r-��wa [�Of9�����wN5���vg��C�}h��i�����
?��;�I�6��S\y��
fǿ��$��٬\'[�,>e?@��ƣ?v������	i-����6�Prכ`����f�ݜ2'։���l�!�*
/d��'���ü�*����o4)�vQy�+C��)ߡ��TV!�yҊ#񊆖2��g=��̚��٥�	��N�mj�}S�� |�F� �G��n�_��0h6v7n� ��=4-?�\���������!�]K��Y|�hK��ڱXo��}oBr)5���ƪt�y6�&��et��!X�Bb�aB�?}�����~Ո����k�7^��t��ƲF��K�7Ȁ����fEF��ü0-�!��f�8.���GT��y�$U��Z�3����	�?'��4��q�P�2��̬�jtG�Q�f+c�gt8b���*H-�t���:�7���� נ!t���04��iĵL�b�s=!�@i���ŗ������>�/񆀝?,:p�l��49����Q�Ox`���;��MzR��HP�q~�����ּ��>n
d����š�N�1�v���V�2�ޱ1�`�(>[��Є��Npth��̈́X��8zTC���H���:��A�U��p����UR{�K֘�J���o���s���}��c�p���6r��b��3:�κ"cYO�W<�(�L��;��l���p��o����l�$��	W�\��l|�!ܩd?�pK����
�&=��P�-�� �>�+��Y����� hS�쀩�_�:�_�CrH�n����=��T_����Y�/ޛd��U�O�X9%�o�]f��j�*�ņBv�F�0�ԧ��R`�q�ޖ��`߲	�J(#
[�%�_�<����I�Y��g9�-�ߌ2Z�
BU1��hX��D��3�@δ�r�-�UK��ENX��0�Id���H=��4R�Md���k�z�>������->%��OX	7Z��˘
��jCH�խ��OG����d.bO�,⣢A+�v�9��������~���C%�����~-��D�T*�+��߸3f��K!�s�p��3�a8�d���mg�<�~H���Jan�R���B����f7�eL}8��k��8O $P�>Ռ�A��#sH���1N��'vK��ӣl��g(�Ω�Q�:�z�g�%6�@��'�^�_���Ϭڈ�M��~�
��߲��!��A�F������q��r�盆F�;�������(��ƒ���28��
~t�rĞ�Me�qE ��U�p�s��a)��jԓզe5¾ g�!�N�������_ٲ�݉:X3�?�a��V����5���l��.��.���c��7����a��������c�������-��; IFL�`L�Ӆ �[�]��jG��AL��C�������A��Sn�k�j��~ϐ��Hl'�����ֿ�{
�:�[j\g�fHDcfn�_�ڴr��|��yOihً���f^��&q��\B�J�~f������s�KV�e���:�>�$��i�_��j=Wr����s��Zr�g�U}�y��0�Ya$v��nw��F����Y2�Z$=!dyJ0��=Pk��p�d	����{|Ӛ�z��@A���~#,���EP���rR�=��N�E{�N��jH�N�;�LC��{b��^ӣ���~g� �)#���A����䐱C�G�EnN�?�n�q�2ع e E���*}�!�a`�;eņ4�	�Lj�2�_9rǸ>�y�XX���I�:�` P�[���grea
����!����s
�W	��Ѹke*�Ϭs�u_�7Q��������64#��Uշ�Dt-�p��M�ټ�@��\k��50j��
��l��1��c�ֹ]&�ES��x�.#w�
W<YQ{$�����Ƥg>�`��������ެ
O"2��|�%�fb��q�� �U�{���z�%t�j틬�0q����1s���9�aZ����ELT��A��:/�B�����A�k�b+���0���'(�)�
��B�-�ʡ�#�^/�'�c;ˬ�Z@����qc����?	Sߎ�f�# �b�0鏅��Ÿ�kZ��G�P��3���˙@f4���@�09�� <&�m��S�N4ƃ�+���}�V��Cd0Ea�$wVq%d���tD�ѳBH����)*�H��e_z�-s�`	F�=�9	��7[*)wx_�=:��������P5L��Ty\_�C`Y��dIQ�emn����Ä��0�/�/�
Ku�D��=�����1z{.
�Kt׃�㮳�vN[!,G�yˆ�*���oS|�j�\@�1�wY� M�g���qyM�7��j���K�\r�́�n'VY�1�@����������*n��Y�f�x���P~�%�$ż���DJ�/O�1�^�I�ǜk/{��-�ÜE��Gf:\�i��M�������؇��$���?�|�w*�Q9���v1\���S2�6�G@za�
h5~6����d+�K,�·��m�ue��Tr���>���c@^	�j���
H���^+N_�E���B["3�-�.t͜��s�-���̧������~�e�'�_�=��{�U��g��s��Ѷ�������Rm���^V5X��MwI~,���B"_�
���<�O���d��T��S5os��9�͹�|�ٌ!��	nS��Z�g͡r���L��s���>��1�? t�����JP��Yx�I�ؐ.�$�i�1|[�~N:�|R�̰�C�o𮼃��r����U�]����SԹaӲiI��0(Y�I���I�xM��k��AX��B�8w�:�P�!���m���&1�g�2������&��'���$N�q��4_�4��mH��b[k}���`�a ~vW��ML�ďmX��O>&�.M�rV���"?8-55��9�����Dg�o^XY��wL���j#�m�I��r��ei��e��$��P��%�i������t`�]9�!��>N1�����;�	@_#��Z�S��3����/%g�]�76~�mH֯J�ͨn�
�A)J�?���K;�.�/�+P�YseА}f�7~Iu�FF���sM���6��6���/��s_J%��*���JͰ(~7�����ݦ�KYA�ν���jfg�m�&�׿1��g��$���1������v���0vD�$9"��xPtp�T�Ю���R�(d e1�{ZE����&/@P�Шs�
g���5�G��3��j��VA��"Ĕ��7�����
��h��m]r��
���8{+}��Kǥq|�P>�5Q�j\�oxg���~)����H��$�*����L�?��<踫��2<.�2�HZ��Eȧ� c��oKOQ�����6���,snq��i��,6��LB@��5Z�`dh���oC�`B�����p�ar�6E�ۋW$���a�^��3s���ҜS�5��{d�CǾ�v�bq�f���e5�����b� �VW��\��3�������]�'���m����Dq�1�~X�3���� �Q�����%5u,��'��p�B'�\��ҥU1w)L��B+�2rL��'��z񷁻8Ƽ�S���4���tpaUe3 �|��~c�0!�����Xna���N�^d7�)��YߘɅ!��S��`��ШԿ�E>$�n�O���mGmM�4w���N2;�X����W+{64�8���䦲��-�r��� $���x�4�laH�FW�7b��'D���s�0��g����s��=��� н�6L��
��	 �:��r�%	�2��رA� �Y�:�Gg��x&�Q�<Q��vxX�ȿm|������H�FKZ�1S���N:A�8�H^�-G'�kDHaxivq�Bm��[)>��Z �2��t��G�nK��J-L�.�z�/�7g��s��B�S��,�W]�[^��.
-�t�ӵ��>ʨ��!)1%�;�o���!F��[wu�<�B�y��^K�X���J����P^#6��7H߃{���?�+���E�垫�]�,Ow��\���n��(�,�\P��n���}���s�sВ��/�ث�/䠙�G��+�"��$����oח���$�s��V�v:�$��x3|�v�3"��v��@GLj����:0p����S�w�lA��@i�y6q�1M.�$�|�a����x($�k[z�&d[ۃ9q��.�V��xw��v��E$��/NT[��V̀+ȝ͙�L,��ݦ�wbXS�'gf��rE�Ca�>��vbr��>��b�k�RV#��Dئ�Ѝ�ݪL���(X����6��Iջa���u�x�S���k�'�*C��3�3�T%��U�����'V������(��0�]��f����΀U��#`9<#zS;?W^�yP�QF���<kMG>�zV�]��nw��_.��z�����Q8�����X���}{�H� �1%�[{�p+��0�_NrSq���U8�.E�*L��]+�qJ�Ң-��#��;�JV��@S�%O�ʻm��k�)�$����"Ķ��$[U*Qm��U�Z��"tJB�H���c��Z�=���Hà�8���<�u#��~���~(�|�����),r�:�=%4�5�F~���"�Ũ���P�r�iq�[��`@Qőr�o��J� o����Ҥ���_�Wf$���*8�[Ė%MMК����m��?������9�M��'h��#���pfZ��%k�Vn�a�G}ʲ�3��"���z3�~~H6:Pv�Z0�3����H,�д�|�&�=}}T����!�A��kб´�%g���Uom�Z��W=Y�a��c[�xTR���V��w�~���fm�&�p�����n"�������@��2-�F���_O!���J�[��`�Mj/ �^�W�������=�	����v�oq!-G�ݗV7�9�h9T��y�9Uٵy�!L��L����#QV�,ceS�V�}�~$���]�z&
��R"V��gb���l~�3�hv;�z��5w�o�e�ҿ��1-�<'�?����t�ݪ,��*x���Q�Z���1�Kpjÿ`H漂�+eeW�#�rC��+�ĤYi� ���S$�=��W���;���
i�ϑH}6�E��>h$b�w^ۈ�gg<�PR�m)BKo��?9���1�-�9.��A���MQm��M��x:;��ib���ͳ$�R�	�X}��Ԕw�M���*�;�=�;��� �Њ�ڊ	[y{h �*w���i\	�(U�hX�&s��b�Yn��$�0�'U�,j�뿈��`�,2Im)��ƈ����&є{���%��5Y)����E� ц��Lɵ�!2$3����M�W�A�;�x�fG��#��8��^�e�/�~��~��&���r�1��+���T�ѭ#��mm�q�Fb-A�MDҢ��������9�ߙm4���"Ϻ��# ��Ru�E�0����O!�%5ǵ5���ZiV�*ň���Ji�/����Gz� �Q:��۷W�̈66'�������hZN�l8b�m#(�f���O� ��\0�����w���4qVۈZ�&�/Pl�6h�F�|��U`�'�&��h��Vs�U�������H�_�66����1&���D7�ma��8(��'Am����`�|��L`����ᜪZ�؈�m��֖I�d�r���!��`���u��WҐ����x�E��$R���p�4�$��dKl���m�\]jO�5��^Y�$%�!�?���3[�B�v�r�֪0ls�N˥r����Dp<����Fù`큒�F���+��8R�S�0W*,ah����-bN?�龥M��h욢��7j}�(���wv5�^1��$ x�PK�y�E����vX3�l������,�%� DY�;ąj��Gߢi��X�O�[Ғ�[�U��T�KX���5�x��s���wf&کh���-�^[�EY�ϟ���w��H��ȓe���=�|��
c8	��^[n���,�#�e�"�s�-1,L��;I�M��ͭ$���b"ZAQ�"ʤY���U�N�G����-h��3�F|�J�l�*��Iq�$!��4B�Z~�Vp���nƴ��
�z�N��UԨ�3��T�LHq��ʈjW i�GX�����$?�'�V���{�S r�C-;[���+3J-G���7����#�.F3\��c�6]��ӥU�"��C{�G�U�����ch損�׊��3������-[���0z�a<�=�x9C����"|�ȼ���]�n����)²d���$I�HbT՟\�칔Uo	A��̳<��0Aq"��D�o��~�5� \�Ÿ��Z��6T�����羆jp�旅��Iڴc܆���Ί�+�lfب�Mjm��DOz�n�6[���hmdI���=�֤�䌻+�3k�?��v��pr�����+=��k�،!ѓ�|��B�-� l�F���[���(\a5��n��^;�I�*1�,5�ܱ�/���2Ȇ(6�W��j�ˎ/���ҵ��:1�Ck������l�w6�s�g=Uϸ⡇gL��&&�f힮$��~�>����@9��J�D�H��������`M��*�+u�'߬�WX �%�3)=o�*"���'0�$�q̿��$���u����'}�!�����&��z���C���/��
�O?��?^�p��ɕ9r��S�8(*H�� ���|2Կ�}^���	�(Q�H;�R�BGZ�ù���hD,q��T1�S{�{�-h�=2�"j���F�J�t�ƿ�����Tv^���m�Quf1j�/>����YGN�}��zw�|�m_w�����@���q��I�qF ��'z���HǴp�"��H��O��B�1{�!�oX��`��k�C��v�8^Jpa��vs;�q�!󖄡�#����S�� �����!�, v�.�'�R�}Md���Lm$�F!'�Q ����j���
�z��2D�ȏ�n��Ӣ�m����ȩ�Jr��;;8��Mh�n@�%v����N�]��' ��9C���mb�q��o�t�h3v�=�.7K�?��5�U٬+G�O!y���P����2���V�!
��?�)fVQ�pÚL'
��}�x�6"��\�,��+!��9�+�|���Qe���X?m����Ϛ0�T�"��JGd��5�k���k�gD8�����{�$�3t4K�	����ؠ_��F��y '������_����3i�x����Rg$����{��oo��ˁ�˒��.�@����X���K��^��\�]V�=��ȫG��\Wj��_�k���RS#������H{�/X�"�i���a\��.$��|��0Kj �L���~�-�ЇLRY?=�X�}p�,� ���Gxwd��|a�$g��I���J٬��@�Gʦ���ė���Fi�5ZA�J��@��ܞ�Vȴ��VFL��Zy�6 9���}u�-���5߁����P5��T_%�;=���,y�?8R�Dc!w��1���~L�H�d\	�D6&-�K��zj����_ �,&�X{.��,�Ď@vZU�;�.�j��t��~��dᦁq"�m��_1u�4���Y�����/���n��h�ߓp�(~���w��v��rg�,��F�K4��#`����=4o'
��X^��c�eh��L�E��q(����UT��PVx��˶!�MsZ0�Z��n-� ���|��[�-i�B�2�3�����J���ڂQ���������l���2�~�$M`R�b�A�}z%%6�uv�����џ@�=8�1
Z-n-�Jm���m�+��NF_DKv��֬@HUk�`6�g�ԟ`���������2�aU�bU��ki�؄�$��3r;�x8!� 1�em��N>!3����0J!%s��uY�2������Y�n7X
�M�tw_�"�y<
���(k߲���+и+L=�3	U�ކ(KZ}U�����V��J�}�d�D\���U��= �>^��Ô�;e��!@:�\ukjm�I���v��d��7�Ģ%g��Pk������7�:͍@��_�p�����v�F����y�;:�^U
Y_�,��~��3b�~�T*��̒bt���U�@Ū@IT6ɜU�|��:)N����[������σ�V���F�:	�&h��V�K��=�2xP�x~h��'��dp��b��G�vr�z#�����SۅA�Bŗadא#����+���{b����rv;���'X�}��o{��E��7�$�"��Ɗ���q�׫��c�+^��|T#����(d��ѓQS,i�8��-��OJ`�����pW��ŮM�#MK��P�VX���s@�B�6䭵 ����_����|���[�$''d�-� G� -.����G� ���� �ʳ$24��_�Q�pX��c5�N��a�c5܈��_(�F�>n9ܤ�c�
����FǏ���Ӽ�^���}�|���y��[/_�29�O��$��o/�����m�Y���C7�$����9R�h��<+�>���~����4z�c�5#�ޑ�m?�Y����z��i6�ߴ$���-���3Xz��r�dd%,Ǉ����'���������vD���.�Z�hWuلg���0��o������Mq�Za]�?�yc9��k�rK��Mm�G���b	��l����\���l��l�U����7�Wr����(�SU�`��<r�y���/K����5�h�.�/ff��bĨڢ7�<���Q�@�6E����f�ȳK�"�0���f?�\���7]4����rX���JC�f��z�a|����9\� -�����R��9ߊ|]�M�l�v�D�C��N=NUB���<�DG�`Ǜ�s��H:z�2By���Q��҃�p~�+9�;3�[��ɢ���]=���I��-�x�8"1����o�ɛ�ؿ�~ɧ��%]�0�����ؚخ�_���%������P���PW���hƪ.iR!C�?mS����U��dئt�%�¦כ�c�	ǲ)��`�)�ft��&��UԤ���[�:&��8��p�	G�RR�NQ���.O� �ňİ	^�)��x�9�տ�7GȲ|=q��Σ{l�?ߋ�P?�~Zy����D�yW>�%S�߈3H0ݦy>�r�,qna���L��o���K���g�$ݘ_o�����Y86s3�W�̀�ǫ+�ON
@�o{��)^�D�/���;Z:~c<�[�\�3m�ݦ�����ً�r���Z�w\آ@��H�G��>́X�_p��a�X��羅󆖌`�l���ֱS_4f�ޮp�������'��j��i�F���y_{����1W��E}�%�r�5N�s������Ʃ��?��x�P?�~���C�t6��+��m궳��5�.�~5�є9SR��.ǌJ<�0��{۾��Ӕ�+�X��.G�>;��V4vT���+@�gL�*ϛ`��������7eC3U��=b����k���~��/	�_;�1,?1�(����6#�.U�v����W-N�X�V��k��xy�?5W��~s�~m�9����Ei��~�D�V�I�?��m��saf���(��#w�B�v�LK��|���8��UTL��k"�iރ��P�w�������T0�	�1��G�JFxb�)����o;�[}rd�ޢ�H��~�)2��/�?��i��Aq��W�١��C�{)c`��������ץ���������!�Y�ȯ�Oh{M�����*��n�8��'���xg�H_I�ȈP~�_[(�׮.G����ZǶs��Dψ.^Tp��S�U}ԭ�-k!\}��J����[ژFy>dn~��/�+�������p!�.��>n���ӓM�����h�O�W+�
z��M�~�em�d���f��ی���d+q�ɧ�[8ˇﻄ6K��P��7�p��i��l����F��6��ԕ���y��Ŏb����?:[~A�V�2#'?��W��k4ص��QZ���]�h�?��
>�ox>��l��-S�G%T}���ٰT��Ѱ��ی�=g����N�y�g��M�َ6�e'���ǰ�G����δz�J�zW��ޭ<����(|�6�-܌`ö�o������]�y��ٮ�@��M��,5͛�L�������/�]�������l��[#dC���O��Wg�P8��~G(�����Pq��[J#�|�c�if�ٲ���y6�U����Y�o���W�6��ƛ^ ��N�Ʊ���O��=˃
[�-�Gz�DU�'o��m�����q�f��횫6��w��!6������L��n[����0�җW�t8��B�?�l�6R>]�ӂk��`TNX���G���Tg[dr��*�?��y��xU���z���5�^�����_�dO������ĕLe��>̊x�yâH��t���=z�)�;��o�T9v����7.�Ai�~�)��\I�~�����|^=�=��l��yMZBG�kr&2��oz��A^�_�^�7r��z���װF�y�0?A�1Yɰ
�1y� �3�bv(8�I��d���\\�ͬe?����TF��a3���.�A��&1�
m�����P�U��/�ӉV�D�O����R�g�Lv��F5���=�i#�Ed��s�Ea \	�����[4��X��G���T��pБ2�)@�|�2��S$��6 ��wI���E�v����I�
!������n�����߃wX�Tt���U�-��]!�(��Ě5%�/�v�J)R�S��gPשQ��FA*|��!��(`9��=�.v�vh�xM�XoVx���34��-h̦����ǎ�	��4�~u춇ƌP�%d��������3{_n��t�M�ă(Y�e���x˗h�j���M`�o�h�ss͹>��PaR�)w������qN����Vg�4�Lt�(���s��=�y�{ �x��,\zlŹ�ٗXo!�T���k��F��jZ���,h�<_Y�Klz���P�|�o��GlU:{��-W���P�I���r;;�M���j/�"2����*eo��٥��(å�c�%;�h�5:�(Y�8�Ő�ښQ3{�~�����5�4	����I���a���Äw0���g�;�&��NƄ��=�z7�n����M�&�հ�>��T�O�-@r>}��{�ы�촡�w�5x�JcU»��ln8Ě_䀭4}���5<����=Ĕoa��w�ң�H����~u 巫�?Dw���P��e�%�����ONyﳕr�Q���YY�96�3��`��%je��OM��^j��<B���D����q��LS��5�5H3�n"�����F�*?�KU��l�P��eM�"y+������G~��</?em2peU?Mf�ZEs�8r<*�u�z����<�� p���h[(���ϟy�%+!�㢇|�����<)=����ss�&@�����E[��`W]�����ro�+��H9������a=U���(l����'.��۸9��e����o>yB0(t��L�����+���U�����*��␍�
/U�1�E{����h��wBygT�MU����@��~���bM:������z������c�a��Ѹ����n�T �\ny��Sh]���'��)z��n�F�s��8���^�eg���v
]1E�yd|n�m<2��T�f��������1HB;ꊐ(��#Ӝ������c�������N�-g��n췼9BN*�#?�7A��������R=hE3�C��:�ˑԊ�&˪@��p��/��0��htyJ�#�˹�v
i#8[�xs`ҍJpO�OD�A�r�aF��S�Q�X��ks����:�`a�Z-��G�;_J�!�|���R�vNi��rӄ�~l��L��4�$�5T	�ԅ�1��%��6pb}UF���Ȭ��������� x9 C����<�a����]�^-ݜjr'�Ǚ�w��9z@�@.>v1�4�,'��K��h�L�i@�\ S5�� ����p�i�6��@�E�]q�Y'���XrO����b�����I����./�8[o4�s���w��<�LG'�Q� �H�<��xPprQ��DJw�	>9��۹R!-;�$ h�l�ǿ�w̢qz�;dYJ�Û�������C}yHdʯ�6�/��/�|�w"�lC��u7M���^�!Q�o+�l���B�e�P?�ʺ"DS��x8)�$��mǳ@Ea ��
d8Ȳ���8e�� g���zrɂF�<U<ւ����D!��w|7��L��x=5D�^��F�m2�@ǂZ�6������}* ѕ�5u��_��}4\�����#Z5���F[��/�ʼ�ܽ`ȍ��FS1gl)ȝ�ʛ[@\e�[V�(ڠ��hZ�@�t��i��@&ai;yS�dd�� ��NY�(��к[�xW��c�s��3:��H���]���_{kV֌��"�~vf�%��Ȁ��ۻ���\�_�p�w��5;�t��^�����G�}�� u'�z
s3�h�?,M���)-�T��Yg�P���֝�E�`C�`8��"Ѷ	i8�;:�L�*�y�UtGKp������H�џ8�4.�x
+�B�Jo�<Ў��S��b�GK~h>)%�V��o�i���)�گ��"�,�Fғ<�~���hH눭�·$FD���
��QG@�gX��,�a2<����(��R���b�*��"�Fh��:Қi@��	E���ޗn(�K�v�kI�]2a�� @h��xz�EӷYq�������ݔK��.�~Z*���x��iqq��(�F�������d
o��.*Q��8��>�f�� <#���a䉥�֗Vx�LG��L����]����>ǻ�R+��˗�]$.��?�N,Y��r~{�^�5�zi��`\ݐ?k.�p˿!�����o.^v���9�,�^\�7�r��2�C��f���{�"R	�Er�C�^�������'A��9#�Ղ����E�P�d��� �c���5!��rs~���?�<��P	�s�Qj�(��o�g��l�j2�<�q�X�'Q�<�~h4��-_Dx��fad���(��[D5����X_�������}tr�k��Ú��\��0y��k8�S�s�`d�?����P7�Ե�7᪸ \����Q\�*��WPF��S
W�ъ��G%��8նk��o?B/�1�3�����V��_P��a�ek�J�j��j��a�y� �Ϛ�A&=�׏b�l��TJ�
��0�q[�q����-�w4ԯ��J,$ �z������"��c�Va�Dmb�ƾ���*n(�w��!�'�Ќ�z*����%/��2�G&["�;�0 �������G+�
T<�ǢD�_�Z��兠�Y�' �z#C�Aɒ{��i�T�
�
X���T���a F����ź�TWm�DLE0��ɶᇂX�ĉ�L��w�=C���햇�-�?HԔKb���E$�~;��r��i�GAG*��԰S�'��F+���	���q�\�Qa��a��4�2�;٩�d~F����n��/Ka�@rj��/����eX�5��"��y�S	C�N�Y�S��a�����U���F+����Z'�8#Y�cn������?����������Ř������d��R{U`^�{g�%�l\q�fM�7�v��Se�V�R�3d1��}H��
���S��T�$IÀ���<��-ȦG�)&E� �H�Sn=�Է���J�dŹ��8�Q���|���F-L�z��m聉r+&y}~������p�n��iL�@B�S5$g�˳4�����nxS\�_���.�s/�h&Ҝ�Zp��B�e��U�T���VU��`�=H���������g��|88�]w0�Z�����8"���jx�4L	e^Q8#�WɠFI����R�}�wJ���2-����!�.��a��x+o�����oE^ϋ�k\���Pha��*+��Ȇ��7%>E��wZ|`<)�쎮Ϙ��Br~�l���`���4L��+��+�0ɪx�]��#.c�{zZn �����퐃�4S�Q�\���=��U�(��:<:e����y��۠|Ex-�FIy˔K+��H)�t��Pi@�p�_N)�F�ބ��H��`;Q��Y�0*Y��,h���<a���ŕL���5)E�v}E�T�l+^���+�Р�7Tܹe�70�Il�bAĒ�&g}�}�K+j�j��#l,��069b�)*�>}��=����D�Q���u:�7|w��]�.����tk�N��K��hH�����wZy	�Lɶ��P��Vx��\�kڷ�+ɰ)dݧG�U\$-\l��n���$-^��j!�r�5W7�N�g���r'l���鳽���8.��`���\rp;�}�f�#������J.��/Q�����:_��ͻI$f��Y�Tx���*u?zl����f��X�Hd��wٌ��Al�Pr�A~+�ū
����k�}�.
8u
�"X��z�T}KS�^����fF��3|F��ɡ�/���2��p�O�V�`�w~�fK���o9�^���P*�e���|Z�kǅ#x���.ym�0��w� ��U;�0:BL�WӣrYG���w�bHQ�/��+�zNᳺ�
w&��G�	�l
ts�ۀ�����h��0w��$�4�)������VTcKS2[t�����r�>��i���U�i���=�x]�l
�L�殖��<�R���RA��/$�}`��`��uZ �9�"��Y7Ƽ{	�q�2ږM�G�|�!s$5�5�%`4�V05SbqG���l��:p��+�s���+X	��,����ϩ�fz�!�Q�_!g+@�(��J�Dn�w՜$)�j�z�	k�-4�tf�5� z�/ƚdp��t��(�;��HjfI�dx��"ڻ}�s�\�]>ұH˰
J�/V˓�Zt*��{16�i�6z3<����KZGJ����L6� �u`���Xr1���5d=�W�-38�>S�C�Y.�{��Z�`fJ�Wpq˒����A�%�P߷G7��+�{����lS]Ǌ_x�F�8��S=K&Roz������/M��btڸZ��xO�ȉ B�$�Ƕ�Y��S��W8i���`�_%Wmֽ����=Y�p����`���z�M<w��ڵyR�-P~9�*]�Ɉq���~�p�^�E:>�.dpy=¤�BpɊx!+o��6�X� �:���CLr���`��v�'�\��J�<a���B�r��7��F�4��k���=�P�[��8�����U#K�_�o{8$yS`��9�7�&?��֯.ld g�N��7�W�_����1P��]��o��L�#�E�'� ��KaK_G�m��s}U����@�I7:]~0�d[��F����{v(l2aS� ɿ0n�<�`��+��+���SY� �������銛����`�)�/6sS2<���"�27��6$����e���MY��Z$�½��V�b�{+�����@����7����үf۔|��>߸�L��7�"'���mn�f^��؂Ӣ��u[%�D�5E	�o��e�K�Q�p�i%���F��,�*E�oZ��N|&sd�!Mm�Z��z��sKj=�|�uV�NA�ixܴo��{�m��@
)���_��N��4[+ɣ�tΉ��l�mǫ7�����>L*|����ɉs��qy�S��$����B���K"%^�fg��r�X?��[t�H����g Q�}o퇕�j��/@�k��^O}����MтJ�{\�Q�o���50maٲE�������4`�ˍƵ�Ao#����|�>
l*�O�ў��$R�ӱ�Ì�cm��r�r~:���ϰY��Q˪��H�a_�kSX��h	��3;OښK�
�ڜ�����x��e��e�����L�����$Xr�T�Ȳ���	��l�G�^ �.��i�6�}+_j��K����:��g?�[_�g��e{c�9�:w�g�.O�S������o���N������i�_�Ry��<}]K��o5�ݗ���t8��.��g�	?G5v��Mߡ������jm�%n�7�u)��3CE}�a�f@�?ob��ף_�6 5g�]Q��B�O>>�w1S[�y�~���YT|'���V0�i2�����o#����8��vc`/���y��I��ଁ�HiM���>%OT��\b28�KεϦ5g�\�vJ_`�c�N	p�(|�y��&E�����I"jo,Xl�o���;��Y]#��b�����3erB�?3�Eȕ��2�N��;��������Ǳ����+pX)-��8�� }� �O١����Rx�&���W�3r"�������n����R�����m
���H���Q��T�]����>��@��L]�16��`��u����Ӻ���r:��r�<����#BsN���,f�2gwc�����޹�"x�1s��f ��JC����:�x��h�>��I)JJ}��D�v6n��T��;>>G���N7/�v滸o 2��i"~����K�{r7�
7���&������ty��-_�?���K�<�zr��{�}��L{Q3��o�����)E�N$�X�^|�*�t�H��S��u��[��� ���f�:�fb�T]~�i�� ��%��@�� ���V�f���t����08Ŏ�'Oo�?z�q�#pe�@���o����<c���C��%ܨ������u�0dt��R�V�>Nf��c��{/�A<�Pw%��p���2��w�I��?���U�{��D�S�W��T��=��{yg�������O�ڜ�I��z���.�	���������Y��>�^��+�Oy:b���� ���o��'��ss��jQ��#�"�9]o��nv	�F9E~�������^���	0'u��#
�7՚��A�T���/S�)����Dd1/oʁp��{+`�R���;NmkY���&K���T]wX��^4�QD�H�!(H� �h�TA� WiҋR��#(�A�4QP���U"�IH�}3��%��y��Μ���3�;�Ԭ�z`q�Ƿ�d�j�/��b�D]��|���ߠ�9*���rr&�|5�S��Ai��}Eeٮ�4s޴��íQ��ޑr]�"v�x��<�����U���+��g}�*�����uE��/ܾC�������P���<�Չ�09�2~��'fDDGA.�3B�jL%/ ���_�M�v\���C鼖���h�IB�I�x%luwV��e4"km�|ڙ3x�������\�����\k?O$(��#�t^ԭ�h�-��v�7��zo��|c7�A4��X�e<�x�6���A��鍇}��)�[#`)OD�QM���)�^�b��M/�����?�9���-�K1i����Φ$���!h2~�:4F�pw.>N��^X�o ��T�H�dp��(Ĭ���O�8�
�/� ����E�W$������J���bd���A�V�Iԕ� j�����O��+��W�b�����65C}�Цo_�%�u 0;$-y�������۹`KA'�d4X2܀I<G������E�� x���%܁_6�rf-.��;��{~%�~#�P�}�%dZ����Wz�{�����L�9P� 2?ɲpY�,�Y=!��o��:B4���rvMHFE!߸�K�����q�0�K��䉃�}ˮ���@�E�!hO��R�v��B|�İ�j%���ˣ�s�R�&��2��fv�Z���=������"�0K K���)r��0�������McR�&=�����O��)7��!~)>zѲ��xi���d�7%^�J����}=Xw��6��(x���@���r��Jh�ٍ<��rQ�N�(�NA 0□e�Zg�<�|DyS9��+4[o {%Τ�*S�߫΀�n��,�Ҭ���|=� ?�k��y�$��3� �����J�s�)��b�o<��fJ���9����!�
b���^	V���ܮKhڤ��v��Xzg����t�~���gt��rXO�[?�{|Ů�Ó�c��ϯSdM�[pS����֙��z��W	���s���@(�T��ڸ�C۠�	�e�0������D���DW!N�
@P{�E��X]��������,��b������E��_A������	�׳	{� ��Vπ��DJ�66�f���Ok�^��N�zǷ^I��q�y����&�����F+��� ˽�騙�q6�Ͽ�����s�2�&
[%&-ï�.(�����������T8w�zM�d�~�I�A��qưbjV�˶�OS��[/i��*���ɢ�K���Z|%�W0�-�
�/U�b$ҸI�c#2�-薶^���SG��h(-�������pU�h������e��<V�E�<u-���n�P��ҩ�k��haHx�S1D��8�rOǁa�v�<s�C'�>���>_�y!H�DCH@/��؈3�+�z�Տ�(�HuvK�<jT21��J�'X0�ݪ����,5�B���j��PB �(q�;SY%�f�������^���$Q�����ձ���\�)�'���jk(��t��t'l뗠��}vQ6V�zaݚ�C�eg ���P�
�Ż�՟-��n?�]���Yz�j�NT'��<n<��C�e^L$S�_����X$;u��J�ѷ��-��h�n�~���sHaIT�ț�U?�!����`<K�Rr�1�ff\ ��Iߠ#0G�?F���#���>]�;�t��.9����0%7�1���?��"�F��g�����-�n{��tp<�/�0���qm����!�R���rT.K@5�<m� H���+뱃	�9��W�,5?�ZH�$
]�k줷u`���_�W�l�Bse�Ԩ9�+�7Ⱥ�$�>JW�o��_�Ʉo���RwW�+�6wP�'C6���3>���m3���Jw~��������P���ԡ�3i	E/��d���s|6����U�w0g���Y��K�j�˄X̢���(;@r�Z��rWȢ�q6�� V��ʻ\;C�!H]UC�b�GB��ɵz�e��Mg8K�[������0f�s�����H�j��j�!������2�|Syʪ�g�\�Fi���Ct�]��lH-��E�FC����o)N�����Ы�U���ڥ3l3C_�xΕu�-u�}����*\��z�؟����4�v�t�2h($���U�Kg�Fw�Ja��T,v$�����B���6BCw#{���GGk>͆��n6N��Z��^�Q�� Z�6l�Vǐ��_��E�V\�]TQ�ݵ@�^f�C)�[��|E�5F2�-��M��X����y�ڦ:�����=o��C��0	?МJ��A��[�>�[e����#JD���P*S��]��A?��
r�~1�fae�1SR�oY�`t���B����԰�����I}=�ϸI���l��^��=^��.�0dL��ک�؃������N
��/��6�Gw2<��{P�!��ۻ��T&���N_(��s.�@�X���||:��Ma/"�i5���tt�y��JF������Yv�ث~��'�e$b�8NC��Y��z�	k�fS�W�%�d�Z���j�R7`�T�:٬�A�x(%(u*}{Ii��?����V�K�`�K9�@�W	z���1%/�����˩J���U����L
��-�pz��Ko��Y�����_����t+��W`gU �<Bl����̪u�?�'{��J��~� )�%<iV{��rS�L.uKd�<R�iٍPr��a �מJ{�zx��;�=��x��՚{�3��WKXm������R�0\Ѹdӗ���$2��)�o�Q:����C�7�H�@xv��>+3�#pG ���;_
g#g
�a�D�@k\�3��	�ǞI��/��������(���9lzY����Y1� �U����m=c��b��骻����Ep�=)$�:�?#��z'z8�,*�U���v�k(����X����s2�yz��v D���z�*�HK�rN@K��^[��ל��\���Lsb�u�w�)n��g���j���ʖ�Ѣ�*�qȄ��<�,�B�,�b�
5鷚��s�D� �d�j��1L�)�8KΪ(z�=�P>��UX*Lo�$sx�m���)�`�v3%���vY7�*�
c�r��]ggX�~���^�k$�l�{�tY<tI/�2Z�b�=��J�J��r
���~��(��qL�.�7%�o;!�*�v���(��L�OK�����D�h9��{Is"y+�� �H���~`��֣_A��]ٹ�u-*��V�nX���ʼfr�Nݦ�9�5Cr�u]Q�.�S�����Mx�[�Z��$�{-u3����@�bOU��c;ױ�kr�e���@7�����9+s��h����in�y@��L�P��X�F���mY��>h���g��*�Z���<%�Ώs�'άa켖���oJ�Նv ��}��K��r��;b@����2����}�;?g����F��iMݙԖc�����h��"��-N��ڮp�y�X�EI�e�DRR&	E͍͸w�L��������3Հ�=�Pָ��ꁤ����|��ٜa7nΎ�d�E���gI~H�(�����nw2\/(<DR��"tif�wݙq�P�z��GkQ�s�:
�Q�<��;��aeƵ�'q'z�1�E������H�
����,<bN�ː;
A��E�
�˯׵�e�Zv.�(��	H[�z�Թ{
�͡>!`e7L-�����kĐ��}���8P�$�ЊfG4R����~��Kc)غ�R��Ӭcy"�S�bzz��2�Y2\	�:A�s!n(��}�;y
�li���#$=-��6�6w��ؤ�|�W�wxlSmr�Ô[��]3�f_5qr=��g��,��|�l��	dL���L��:�!O��&7,���j�(��(�U�"^��Sz_+��|�p�u�0�;}��M�m>�[tlk��<�6!9>�ʣ����홯�t˓��������P��K�Z;CIj������'��w���\}�T�q�N~���ǳwF4��Pt����L�4mU�i-ď��^�_�Ѝ�zS�C$�����p���0�S7K�&�(/�x�N��l/A3[�_� mh\�-�����h�d�*����;3�& .�hi�	��j?�Y./ŔIr������|ܱ�e�5���_��3�����Q��T�f�eh
J������c7��@��&�HjBdTp��ՊR|�y3�'P�m�L�mO��;q��bn����Y~v��?�bʻ�V��T�w�t+q�lu���Ro���������&�h�z��d�o�iI��e��NS�'�謠�����v~S��m���ٍ���k�6dڡ��̉�H�c�i�ɵ�`�D�2��|���+�#�^�ve�2�M{����� z޶�jT�vY����tV��I�A���@���ho���YW������ �S�g��c/�8�j�5,�O����y�cPv�{���{>i�A��8�=v1�Jถ�80k�uM'ue#d�(87[Q�:힑��]l�������﵌�UY���p�p��]�C��:B���"=ߙV[�>@��Е_FTB	���w�&'Q��,컩��$��u-d��s1���Tu�M ��fW$����~��	jgG&���Qw2о���h����9�[�Z�ֶp��D�X�J*�1(������\�]{2����]eZ˜�{�ɲw��8iCnւGy��[)�ֱ}.�>p
23���-K�����` �=g�_Wn�	=�\(����)�M������w�Y�!�J�FM��/�&�k��N�1�PJm5�>�_{{n`�|N�
�}D�~�G�=mZ	#wP;sF]����ye����pd1j�u�N�5��w���=���6�2��%8�+�����&�8�I�3����!�3��!�x���IK�#.�IE�ڔ��O�?�}��ǩy��xJ�����F8���4��bN�~e�n&;W��Ƈ�o�� 3P�@�x�D�E�h�v�%:}ss�\��>�x�qG|�D�Fy�p� >��M2��c���]��"7��gͼ��Z�J(�a�r��K����w`�"�=Vm���n2M�!��aa��Y~�ѧ�NgM�ou��l�����:�p�$9���/��x��߭�s�M/pn�Z0�(���h�)�_4�`pj5E�R\��������A�Z��3R��k%~Z���m{qjâ�oƗ�LM�_MI�ˢ�\ ��Y��d _�\[Ϛ/�7�H�2|�[�^�������(��l�"��S���X4�,!!�u#�lnvc�znH)�LgzZ�0|�c�xjBM���� yU�מ��͵���vc��cC�4�C�[��/J��;�K�m$���z�ގ40"Ň�����y�;h�*�Rre;��k��%Ud��္����w�H�i3��mEb�|}���eQ��=H}ф7k6|w��W�i{�q�`���Q��p#&m�+�P�U��8�Z����9�J�UM���Z�M��Hv��)����4�c_1qy�=�M���I��nqw����Q��<�$%��q��ʙ���`�gغM����K���R������:��k��-�����qi%��K�W�;���f�w�xX�2 a����c�&눔��5y�,�B%�J�% ��n�CDt����!��O�O]Y�ܘh�c�7����#<�C���+ F��`]��i�Rmjʥ�0�t,����/�-e[�3���$�M��&h�.\�[�}��5o��_�>�$���p���0]\�3󏺱ՊU�6��S^R�ˉ�m�Կ�0���xi�������-F�9��'EJ�.�tI�� ����ulI.fm$_�T}���	�����@{�Xj=�L��j��; ۠K�!t1����� ~�RQ�b19(L�Τ�7'�<~��ĸ����XLE(�v��L�fP�F
�j�۹���#W/���P�A� �0��!��>qS]�gv�hz8�Q'��4NMX���;08Gk�pe~�����iiT\x��UB-}��[t��S2�B¾]�v��}�h�_f�mod�Y��,'JL� ��쳔��OJ
گ�O|��ږ��9�v�֫�y��i�c6I��{f�*�2�y����_3������'��"Õ�[�~����k���7�ӊ6��8H�3s���pé������ծ�s�鍛�)p�D�&��B��c�u��l�)jo_[�-�٨�Am{z���e4Q�$Ƌ�مOI�i�I�~bEߢ��c�[��Ԏ�%$��[�.ʁr��lZ��}ݟ�93F-Ye�Z�h���2Ӎ�1k�З�� \ZZ��/�C�&�i{��_�{���wK�jhSyX��� ͎�66�ʰ\>Y������N)����^TL�k�c��,��p�3^@v�`2ng�_��(��k�� aaHQKlb�J�2�*�6=mb¬��'�	N���򏿳�.^��3U=4�Y��ݱ�D
rc�m�r"7+�*+�vP�ؾ$��g�!��<��t'�c��mg��l7Pn?@�>���O���`rZ �B�&Lz�p�o9h���H0ifm���E�lw�YrKZ��Dŋ]{FԊg�`DϮ���S��tB=:�Wq�%M[j�q���s2���wG#0����\��$�������@��T׈�̆��|�<YP��a�Z�N� �z���r�l+z�,�|VJ��lQiز�~��O��-X���j
�! ��kfS�z��Ļ����<�ׇs�A;��v;[E(Yo����S���-������[)N�d����-�mn�KßoQJTN3d�2�샶K���q]�A%�����w��)���W:ھ�9�E�����3�h�Y�Ran7�������L=�ׄ�[�H�κ��Μ�g6�Tqī�r���K$>k�H�4�3M�j辩�*����>?A������f�W#����z��.������T��0-�B��ƧQ��2_�>�nWۙ��:v�	OOdR�w��6��~�̮�+�ŷ���5�P��~�K���`�7Q��j�ɑ�]w���6&��P��e�ۼ؎Y���-3��|6SR��;�P����'ބ��K9^%M�R�٬��>��؂���}���W(A%l�֜;+�掅k�t�Ǫ�.q��R7�������:�k���]����������t#�"Q�"tׯ�u����d��.O�����P��Z�`�ijP��wβ���m
WV�n�m9`�s�*B��T�\�V�/gsg�o �t�>�슮Ռ�s�H�_�#��N�������'��p�4�~�ěw�����~οʤ���w?���'���:�y�}u�_����O�n��.ި|&��Z!d��n��ʃ��+T�/�d�f\f\<d�>�|�Ju)it��z夾�-�&��SL���w���A;j���A��xv�a�[?�Ө��L��o�]���ڰ3�n$J*�����d��\��@���8q��Yv�oÃ���ݠ�Z�����Q�a)��>���;�T�������%���;��,����5;h�3�$im�U�V�B Gr�֥��H̹�3�������9�%���Le���ߎ���M��|N��:1Y>�y$C[�����o�у�2����$ILWS�����r<g���f��<��%��!ѐ-����$�[Rɸ�+y�����	��ߚ���t�@����w�P:9h
2�D-���`Mi�8	��ƿy�mO�(M���圻�}��/����s�F������D�!ӍM8�Q�d�`��l'���K�2�ވ��/"������UW�试�x
H�~��yg��f��G'�%%��Ng2쯁4����ҹ�9��!�*�#)�6�Q��B�t��_+���ߞLo��*(�B�O0R�au���=qФӺ(X���Ғ܏�蹀/��*����CV�K?��6j�����F���J@eS�=�S4"�%E�l�+5�b��8h��"ٜ��|����]��%��`$�)��6,���b9���;g���f�?�F8|6J��A'�u��#�Gs^*C��7!���a�뒔I�*�ʏ�U^l���n�ǝ0�t�k���UG�����~�ZG�ӆ�Y~]es��uڬ��L1!��PL��wL`��E�YЙ̼O�ב�����������/˳��0K��3%ph�>��,��ǿV�sΙ��A���V��{�A��# @�)�cl>?r�h5N��8Hm��a�ݏ�'@��Q�m�[���]Wy�#`l0��i��4��M��Mq�F 9z�Hj�j�NÈ��7����MN������9v�K�3m���(��Qg��9f�^G�˦�g�i/��I�Si�Q+����_����(.��k�2H�(����D�y����!����k0�tU�w�}���N%�bs4sÊw�d�˖nAb��+t^93� ���
�<f9ױɬSo��*��w����#
C�����9�����\���� _���j��ր�(��>�%%?��āy�dx�r�b5�HI���V�nʇ��߇lp�0�쟣q_���i��f�i ^T�g��ĝe�X�d���`�y隚�9X�	�����{�hi.O������I��cqb��0PA���°@j4Nr	4����ns�R��Nå�?��g�Y�����m�������\�9�m ��{͞2_EnoY��ra6�S�±uq����P�����d_%��,2�F0ϹL:[�&��Cۤ�/Oe�a�:��r�u��#t;��E��ﴁd�Z�uo�����xi�9X���2�W���!��*�UW�S�o5�B��� Ǻ�G����2 Z\�|`9)B��pd���� N~;��A,��_ י�̆��ll��F��r�y�������!�L�|/��&�vQ���8��.����hnT0ޙ�|����4�5���$sr(^�����o�K�U�BH� X�hin�'ꖧ�:��/�r�Iv��A��$l^�=��"Vt�r��SL\Y壥K]�[����O����s Y�I=ۘ~��[��C%��D�'��NTn���A{�	A�B�Fg�Y$�kˤ��|9k2�&�`qn���<�?���V�H'�����/
�s�'Hk�D��t�l¨�N���6�'�E^U������\M���޸�,k�P������BZEy�-�x��3���B��|�����(�t��*7�&p8(�v�hk<QV��?H�"U9O�3�"l�O��͘J.S�^�(R@(���=%[R����IvB���>�e�����˲tr���c�u�|�����=�������= ���~~L	9��l�� �?gn9�~c�h-y����(�g1븟O�6(�\��Cz��s;������ͩ���Ig�j��BP�&FL�O(���͓M�S`P���e��FSTp�o'�Q�/�5�s9���Y�Y&�)�:o,������aA����wQu����Z�{�t�0��j*{�*2�UQ˩l'�r�s(l�#��i�o,;v�^R-���N�H����y��/#����ED��`NC&o�t��K�y"3\{_���z`�`LJ� �����L���q͉�k�c
x0R� o|�,6�SP]�^��娷�Te��zY.@~�;[N�&�n�j{�D
��No�>b<��F���Hq�\�d�Lq�(�#�m�F6Z]�UU��?މ�a�:ߤ>�eA_���+u���?��A����X�8W��$eJ�dE�W,�lb��9�
���{�l��$oh�l.R��O{x���B`!\��f� y���֨����|G�ޞ�u���#���eWF���O�\�t����<]1L�U�(\[��~E�c�ȇ��-c�E�%����e7>�P�}X.�����\��%���s��T)P6M�V�7"2�B����>/�V��5�Z�W����q9<T��(|^�	_�;gj����YH6m �5����Lf9B�B���|�����,�#�<Y�o'��)����D�3�L��i���(�
����<�����}�>����/9�nb���k77h� ���Qr\���R�-N���©FLK�F��W�����e��1�͢���2H@��$3"��L��̣��x"�tY�e=n�U��T�a��
P3Z�?c���v�L�׀�A� ex��>����$�#��uP���e�{L�cCZ_zȍ�4e�=�A뇃���{��ĥ/�ġխ����0��9�a�,A��=�t�3�k�2��Ƭ8-ۯ@�乾ʫ�@���_�Bc,�{���Qwl�-�r���&q�&�u�Ɲ�K0D(���S�
6�����a1�	�Ɲd���U ��p]�X,�+Tl<Q�|0@o��]�g�29-*�9�)����Z�b. ����E�,lT��2$�v���-C^hS���O�L�Vޒ��q��PQ3ڌD��8KŇ� ���	_���A��T�v�,r��ic#z�vȏY�z;�-�K�~?�6X*���%�Na����ߒ��hsU�P�S\��
6���.³H���4�u����yXlzMV�:�	�t("wI�\����.>���Y�C(h��l�ޑ�H�
�(����7��Ӊ"��K���п�أJ�B��t�}��#7�*g�l��!o�z��P�S����xwJ�,��Z%������_sǪ����$�N�h14b�2qV
>��s#�����Q\�v�XpgD��Ж�}e�]��	nЭuL���Ll)��$�������6�����*�����m�e�����=�5cK��X,+��M�%)!�_���k�%45�;4=tl'�R;t�y~/6>Ȃ�����L�n��}��	:��h(z'�V��c�)�����3�!���q�^�#�1k�~ิ�d����bt�W�1���D+����wN_x��-�c:��$�@�Y?����H�1S�2�TKsπĨ	j�\��؏�"$ſu��F�6x`͖� ��[UU�G�����ȵ>��h�OoLqs� �r_��j�����]5(քa�;�$�S�����*��l+g��m�r-���	�fF�f�Zs�ɢ�C��x�f(yLw<|�_�J��G�����_���Ϡ�&�͸#�^Vmʯ�
��:Pw��a�+t���}|4��,��������(@�_Ӥ��lFt��3D�saI ���-d���U���F^~�ːՋ����(Mz�lW��!��0��:���������^���n����O՛��P���'�lp�%���NH�G7|�a��)a� "u)ZKne�]y����	����(qLN�����~6�u�I~Ui�G����PxBq:��d�6ZKE�9r]��d���ha�tv!y7X�`u�Įz�/��#iePR���+��/�ª�3���ud��\�.�i�>Ѓ�C~9�7:|`�	�/��@����;"h�p.gf�[�*q�A>e:�`��ї�5��N�-�_��l�<��Wu�*6�ax�`����c�a;����W�Z���g�6	�>�Ӥp7�d�:���2:G��ot�8�3,nx=�ڀ����@7����Dn9���� n;�	t�
9�w�h�g�T�'��8��x2^�sB��t�)z�Rԥ�?}a}���%(NŇ[�����i��y�T  �.�H	5W%´%��a�z�&��j1ɹ��TNt��}c!�p�.���:Q(S� /�2l�� ﮯ=��ܾ���AL嗶���S��,�0D�a�u�.4[ �N��ܯIQ���P�, �v��Ƅ�Y�����iԃ`v�"������,��Z������`	�p�8ؑ�m���
�I��}�����Z0.�>_-1W�.ۨ�����?�U��0>�N��2/ҝ��`	m���n���2�I�dx���k"�OZ�f�҃< �/,<�}[t��-@)z�e��*p�d���G�Ώ8l�e��z��� u��;_/�Uѣ�5��ew.�ܷmS�W�u�~u�Jp�<Yd������	��+�x����?�Q?F+�}w0yeb�q���s������.��Zp�,�ʖ�]�B��<d҉���=i�f>Z��M�杗1;M)0Fܠ�rr����Ih��+��W���;�0a�@k�s��v�~���(q!{tx��{�_"/�.���<����"Z��W��[z� r��u������⇊��ڒht<?S�����4������������KlE���� oS3#��E��Wâ�k��
@ւ;l7���<	 ^=��UfiFc>#%���э'����R��wu^(ȋ��)�����֗Z4m�JZ]��=�H �қ�>g�� �l�ڞ(���^/������>����N���$�����z����P����u�[����[txc�`�|CSN<�jE�咾���bt��T,Әw�����.��+
�6�G��Oy����?SO��V`�0k����{s	-�u�F�YP�8c�q�4��� WKޚ~llu���eBh�C#�W}�����������/�<���Og��1�U4|�yTel�����v�w�ț})�&�*�ox��@ű'���$ �h1���'=��;���G#���A��?W�t����W��`es��P�T(Ř�wc�$ Đ�`�C��aq����?	��<��U#6O	����z.������Ur�(�<
4�qZ�����@��[�ƥ�z묪q�ړ0@G#�GS�|�cSw�f�]�l���v� ���zP�]��MSSݿ�&��>��N��n����G8Nu�M,�e�Aڱ�N���ew�vpS�[� ��9�?1�她^ǥ�u�X��S�}VFj�	J�������K��s��j�+u?��/=/N��y�싍 �p;��"]��E;��p�dyu6*����QF����~�����bc�/X ���p��K<Â˥��`k"��Oo<�*�3�L)g��!aS�UU��#b�exu��瀨�{A.(�H���ܻ,�� �2����}ێ6�R�	('*��v:����Q,1�79�d�F]�{�= +���`ݯw`Ƨ��{�%�a�8S��
��'��T�gS�@WM��
�œ���.��G�z� �v���t�d������4=���u��,��evڣ�%��"�{ea�jQ���/�]���/��=�4��^��@'�R��2C]��b���6DI����P�~E��1)��r�h��a�*��<A:�[�lD���Zk�s�ౠa��}dk�[���D��	�7�0�����hϭt`72��]M'(�T���i���D�%�;JT�dqOr�Y�[+�	'�r��_��T���>G�(�~��PC���Pu_jG���'�l;��	���4\\%ܰp�]lA*%�n� H� .��B;���4��>x�0$�Z�k�+jKQq��J��������,�M>��tj?��HH�P�}X�ݻAj���&!�~*���P>����E]��{=��ț����s�|;�q����'�͍��Pz�����,�{�y��j���'�P�`�B	~����M*	��M|��x"�`]".n�n��?�H�ã[^r�z�i�~*F�B/U��U�#��h%�
1y�ׄ�T������D �_���Ǿ�0M�ͨ
�ڳ�}�~��-�9/W������^� ����Y����c1�ͫ�0ǣ��& �x�e��g<���Y�U�c���_����7��֝��an�j���ZGQ�����Z�[&��T�lR���f�¦Uk�M9��Ϸ��OR�����(B�Oۃ����7�%��S�7ٛ�jTF'�TSZb��<%��7�y���[i $�@p�5��c��%��n	�VJ^l��`�/��?rs�D�ǴD�I��
��<�r����z�~$����"����x��|Ʒ������-<���ƉP:�=1��^��4IсmU3��wV5;��z|��$�C^MI�D��w�4�yx�$���09H�rs�|ص`��n
��gnF�
o���� �O$�28���!�������3�] ܯ��n.A��2��2ӄj��E8���������V)�c��2T�%� iVM�7dK�kS��I_��,��($&cg?}"�N�CR�G"��?��1�#��~i����k=�m#'���� x~�#�k�H���H)T�� ��b����Ӄ��ā���:�.����@@�8�9�� �~9�B�K�,ov;�k����O�e�b��%�o���|V����@uf����S�s��	c���b�d�a��A߄q}��@F��7!ҷ�}����R_;����[��~P#��}(j���o�>Ãd�eޞ�9V�v�AS�i��#�e�����74�z�N0 :�����V��S(�g{�z�T���PClݼ�M[l�E9�3�X:�?5UX�]���<��I��Jh� �R
�> �s�������SPA�Z�9vͻ?���'�F!��1��A#>O��N����)�M��~X�]��7P1q!�A�,|+���{�fp3��(rU+���4Im�' ${�S�Dǰ�NFS��=u�:s�K�4i>pn�/Υ ��E�.����W�l���)M��@�4u]��y��?ב�Ù?2q������4Y��TU�ܿ���x��,���b
C/��9�\�L��tpx�!�w8�ݑfmo.�g���&���aO� N��y��#5/<�	i�GHڽ0*���q�%�L�	k�����geی�ay�4�T������$[��߾>x����f�2W�MJZ����Y�p���\���R��9lhj^�_b.|��kH�3�vz@k�?�W�Si'S�-������3�A� �8�6L�M�q|���p!�0a�:���h�#FU�00�(;X9>i��o@��V���b�u��Z�!�|$}��#�l�M����vK!'4q�S SX�3��I_��D}
��E�W\�)�n�h����=�\W�.̑�|��/�������:؟i��� /Uד~��z��X=�l�cW���,�ۯ�0|P}���x�sN��`[��ѵ�C�g�]��w�#�W������Ǹ]�8��y����^�:\�Ҙ����F�X��:5'�����z���4W��� � ������/Y���΀?{��Ĩ��4#8XS��_�k���2^}*��?��L/���e&4%�4�mì� g�*�ڃl\��(�^JP/��y���0�� �{���k����U�T��Eg=�6�o�i3k�"T0>��^?��o�?m)Ef�����((U�/L��i�w�(D(zI��7�	)�+���I��� j]�sW�MV������~c���GH+7��2�@S��0U�a����R��C��G��� �mh�{L����P�@n�#%�-i?{�Ԉ׷��H*m�@�������R�7���!>��}�Op����[r�;9���A��[��d�{�v&n�e_Z�A a4�pE߬�C��'��	t�w���Q�j5��ξ� ��x�yՖ��N5ނ9�?����������B�n�+��N��A����z0-��qROQ�5�*�1�?���?���A�7w�t�Jڟ�q��Qh���@�B[$d��7%BkoL�tA��vF긹,:'@9��f�0�3�}R(���,�鯽�ϋ���TV_;~d�q�z��t�$�j=ko.h�X�Dz��!�ɍ�;�/pC�?�l31�Ӂ��9��2�$���\lI+L؝�G5��G���Px5E)�����#���$-�Aj5��H7�����ܱ�Q
L#�k?���[ُￒ4�J�k@��6Ю'���S)��]�B�}@ZMӢC��b˩3�h
)웖}l�{��;5�yv5r��$M
x�~���&%�^00�م ��(�L�R%���xgi�ފ���m��Z̓�;i)'/%��,+�ݨ�)Ы 2�u@��wo�n0�I-�r�Z�� ����f}����~����H�A�ƶ�%��m�*�#���N �>�l�h�Tl�;AQ�B�ms<��r^IL�f���v�8
:�~�ۄ��������z?�`I"��"��M
���X�ݙ��A��2�mbD$T�wTT��3���b��	�fF/	S%���=H=L�7�tK�m4�޹N�(��@$�Ѕ�ſ��*�ȉ���y����v	���Z�_���N��4B�XJ�X��&�hZ۫e�ua9�#2ə����!�%�,����BH�b��ECjGt���|Ճ�)��m27�� �*!AB-��mz���^-��+����7q�C�C���zˁއ6�n�:Ԙ�=8��\+KK�A"u��9�qɚ��q|]n��2�=�`���c��~�MR�m��;�[��|q���,Pv�jN�Dڟ�ԽW�%�p1�cco��D�yev��9~�5�I�B�3Ld�"��}i-���8�y~�s[�|��v	4�<�]m簒���R�A��=7r��eZ��/��F�U V��'ʮ�?���-7�O	+µU�ڞ@a�3�N��llzn~wJ��m��z��-K���BD�w�?w���tr�1u���,R��À���Ԛ��Ȝ>oY����Ly�� ��&n[l�I%sڤ~��+u����o:@�i3�Y��a �.ͬdE��F9��%���^:��]kr;� �V���w��>��=~OC�7%�BG �a7  �gQ����023d\ϑ�[�q����֕{�պ�S^�:EJ6��/�2��sޮP�3~wF��L_�+(�y4S��@b���k�y��0 �\��[���Y��߶0�&�.���A�V�#�O��������� �8��]��v�l�����P�*���6�'R��6�٭�Q�ɴ6�H'�݀�A�����/G\�:���b���!{�u ���o����I!�dm2)���O K��!�*��A׈�CHo�v+)����&�( 
�Ŷ�/h������g/Oj�;�<9�V�,v����@�=�W�� wn��'&�_�.$%�X�K0T��ɿR��M?���WE7r��r��IG� � 1L~� ��M�\PW��r�D�Jf�1P%3Q��5���0M��΄�U��J�a�Ӓ��M`=��қ1v(�кe9�!i�^�J��[oy�&1���騖��߈at%�ϯ�!��c"J�5&�eT�!�������ހdF��p�3��ʪd�lu���<�п8I�q�����f�� �ӃR@'ld�F�^��'���J��y����f5 =������\�_8
���υ�I8�Vs�;v}U�6ټ�J�&�$�q��<�WL�Y�SF�c�o!���I�����J{ӿϕ�^<�@=�}0:�V�>��5fd2\��KC�1&�ˤ�]����I5Q1� %��$�.g/�-dc�E��nl�ar8�+N^?����7Y4"�!PCk�aN���o47�1^l��1�IWy	j(���V�=�@���m�H��{A�@=s ��j޿7���ӳWF��s����Ea=���t|��V�:^*c%�zd|�2K���M���\�U�&�R�����=�t��ÿ ���/��|��j�=!�g�'�\��o���g����f�߹)����j�~��a��85fh,L �-�D�L�F���iY�G�d�B����5�j��Vɤ�H����xř��0�#�[���gؓ_�Q@���$G}����1����=':��<�K����B�GB��5����2��Ltb4�ѣXRB�Ȉ��&���$G�R�4y�A����k��d�%#�gJ(���<)	���qu.�� �%�݂bW�U���䋓�3�Ž��Ѵ��f�}���B:g���ևwO�ݸ�4�5ğ	��Ls	+�����2	��������]���Ӫxr���ga�1r��D�~<��u��$f7�� E�'�������t7����%�Ϟ�$�){�`̡ct�=���>?h�1���?N #�b�� �]{�?��F`JpC=v*��HF�/��O����!eT�ͦ@Сtfh�2@�T��;
�Ӡ��q�T*~��'O����4��X������e��
��H�z��#�d[۾�MD�U c@��G�f�[\����D���C�O�<��8FS�ȂCj")����0ߤ7|ӓ@�x˼#O�6���͘/��k�����싫򋈑U�[b9�O�>�nm�2R��CU�t1am���W3�3��1��f����?��Ɔ�����n%�%@s2�!�!�vQ����2�`����$m��cv�`A��o�������(U�mT<��	�k6ɲ�Cm؋S��L0�4n�*Ɖw�32���Sw�:�s(ö�P�,Ʊ۔�*�CI�wz7eC�p�&�O�b���ݏ �vbg(.G��O�r��G�n�r�-��7]��x��J�q�����V���gGGa��1����%��^�u���y=������$�[t5p����V����/�ѷ�7��0���l<�u@�t���J����J ,rW��w��o��WMn�F�-�}��yaԹD�S6�k�m��0Hlsܞ�#h�(�M�sDW_�݄��`KO�!���"6��n���ytF����f�Ф�����Y�"�KQ��(?k-��kۇܨ�-�,v>�{ `����˶��U��%��>�Z���x{�����u9>r!1xNs�e���ev/��ǽ�^�K�X�C�9��۰��\�?��: ��k/���R"��H.����J��%( %]��"ݢ K�t*�%�,%� �t�7wC�_�s�=�s��wf(��s�7	���'9�vi�X����H�>�^�H������"1q~Y����yj;�|OFC��!H6�;�`�F|��]A��CbDB�Њ�,ӧ>w�Q�Ts�{u��]�ѺS��ܰ4Y�	��=�1��쏔���L�����c�yi��Yw�ƆR�@'���DP���a|i�~�-�i����1���6X�Y��hN�"R.��Nw≡��U$��oP��M��=ڍ]S�v�#n:WD�+EI�b^7t�Qü#	Ult�l��ԑ�F���c!�5mn����5�Ů�{3� J��������:�i�9��8��#�6̈�L�i�����@�>�Eu�}l`���R	���c��J�k!��aR�{� yB;D�7�	;5�sCͥ?0�ۅ�6�bRo�g��vUT��8��ؔ����r�&cI6@�_��O!���D]�f�
U]�(��f&�nSQ&�W-E����.}���c?�f�p��뭭wd�ˠ�]�%��#Ԇ���Z�Zq���~ƙ�E*�H�YЕ����q|L�߼���uJL��h��PxVK��v8��n�eu�1��:OqI�����a8����lG�i��Q�交5��\N�g6�~B�U,��C����Ǹ�!{�w�=2_��	n!�'sd�T�x��Cp$�*�*q$c�v����qj�� �^H@_mmKt�Z+�|փG~Ş�J��P#�?��qj\F ��̫�O vf�������F�����o��8�0���I ݰQp� D3�=I�W��z#@/ �_��C%��,Ф9\�&m�ՠ�	,�'k�W'�b~�}Pu�<�;0ʔ/���s�D ���t'�u)� =
�Ylm�pd��HB����N〛�W�������Uj�u�y�%����W�X���<&ۥ�VӲ]�;�+�&�Ʉ<�5�L'3g��l��B�Өmr�z&� ��CYmM	��z+�ۛH�yJ�+�����F�x}�J�l�����*w������x��ä������m9T��zik7��ÏA�r��_*A�i^ʪ4o��!�*"O� ֦��x�����1�� �rq3���cs�{r��(�Rq0�P�nlc���wb[�m����D��ʢ����mV�MSl�.�Y�Ì��=���o�ѪK�12���8�k� Z1�fT�|�QD:�m���;����"H6�[�g����`�Q��C��;b�������'�..���� �``��Dx�4�"�H�B�Խ7>ON���7B0vX�ۆ��� }0�Q�zB�ּӮ o[��2�j���)�Ü��q�W�G*��v0@km�MA�שּׁ(~d!�����{R�GI{��8�x�Iu���Z�Y� o6��d�w$�7I�3����/�ɌvMO��?�j�'��a��)�܌��['D�g@$�C��{�8�(��e�-�ݴ����~}Q�� }h����7D��еH"/S-%+$�t��ZL��ag?��p��X|���(k����U-��n5<�񿕌`�a�����RZ��(&�w@��n�ŕ����9P��:p��+9=r��L5K>c�bP���܀բ&/���NO���D\��ӎ��T�P���@�\��˱��I��u.#<[�vu�aܸY ���8!�7��;Z����`���jT�3��b?l]��酏-�������Pf� ��1�^C���c��l3D��2��Ԉ�c��c��f���?<�҉WRs�
�3�w�Cϭl������L',��ޓ�$�p�g�<jl�н��Yr�h�tk��W��RȍIz%���}1a;�?�M�񕥷�����"Nf�&�j�r���%����RWX��3if#�0��mr�?�|F�˥NIdo�μ�X]�u����Ҩڭ��V�f��ٜ��wh�N�1�[uӂ�Y���rE>��K!�2G�Gn��y�Z�]�BN���Fg�;�iEO܌�l��%�*��B�k��LFH���s�`��\�����Nm�ۚ����ZLh��(��'R�bKH�[C)ŭ��]�1hA��JE��6l��%���6�~���f&��dG�.�-���ծt�SO2Xte�$�Ͼ��������pnZwj��,3��e�rKwƻX���PFС����PG3���v(č��?A�k_��5�Ԭ+vtw���7$b}�WuD�}��$�@e�e�ᴔ�:`�bg𴔣X4���MEs�����tQ��>bzz�h&-��V>�@Z/Cd�!~���Z�(:��?�`,��fe�Ed��\=-��z�����l�~�;3:��W�Y�'��>p@92��z��w�Թ�ƚ� j�c�.��i,�`\���(�>�c��J���jT�
8�y �M}��2C�#��9O<C����׮�V��7d�ȡ�T�E[u�9F��ͪ�^���̚�cNL��{<o�$,/Zل��_�-Z>eƻ�J�v���K�m����v'jm$gznѪ�ad��.������뙘bg� Q���>7��gE�E�X���d��k`��ȪC�����YA�Ze-�Et���^?�����w߾��;"�G:�eH�^}�WC��T��3�Lw.t�����JX�w������)�k��F��H��������59�g��~g����T��j-��l~����V��s	~�SK0��9�SɎ�9v��~�G�-ۤ�3��������p��S���|c��$?kRS� FK�.����3�c:���)%Cg��!�ׂn�/C���������T��g�km�u?\�֝�~⸳7u�J��^J�����f��@u�xT�N�����JG�!(�_պ#��NZ��L{I��x�9�#g1�9�!�!��/���\#ߣ�L�:Y!c��F�>r�������=��2Ci-e6&J�$$o�B�l�_8 � ��B�r��?�Y#G��^�|��?��d�i��HIIq��J\�OR�v�<o��U�B���M����&�����%�\Ǜ,�M�B5��+�?v��}���� � UD,�"熜Q�P_��;u�Mգp��X���֐�^��7���R���VMs(��������2!��Uƹ������)<V��y5O]fEr��\�G	���_���Opp����O�f�3?��_+����.-�t�q]��>���`���t���k{{�#�E�d�]U-X��8�b���� ����?H� Z�b5���mJݐ��Rtߤ~��Ӎ�0����.f֧�93�'�	9O�(P]��ΫW��H���(���C��*���y���_U8��#�p�&�ApP{Ng]�`�FpYP���R��v�¹���"yɖ:*<�D�G�ѯ:���4�f��.��:�֝�W�AWz�ZZ�kj�Dɳ�<fh�,EFqX<��Mq<�N �������;�w `Y{�̅b=3��r�]#�%���lh�q	S0�H�.���N�P1�0��,p� �޳o�n��!1��-"�@X P'����!��ZY�Y2+�[�c��CXP�:4�oo�Կ����V{�<�Ŋ��xH�?��ݱ�[6zB:����"qL��r؇�u���W~x�:��T{�9�i����~����>ڷ�����\6���n��dV19��ܝ�\�i�}*H�w��@��cr�2�_\�=;s���<17Mi�O��AH'#��p�rJ���V���1�g"�E�gk�O@�jəו%�����A����<�`�*?:��y�_\���Ä�e���4��}��
�@ꗸ�Y�)(�|���R<;k�F�:�\{�;�ѷ�&ڑ�H�����&�/�<a<��fq��ZD��?m�2�R`S�gR묁DJm�����4�-�S�f�˪2-�
ģ�c�k���	�ڲ�N|m�%-(/s���#��t��A���u�n{�|�̬�}��)*r��x9#��}�2~���������Q�(E�m\��	�[���
����]^�rr�[��g��HgrhǏX�Z�-��������:7+D�G���.;H�%����i�0X���]��eof;�Z��G1���	���;�$v#�6�<�ר�1O���h�)R���j۩:�{�]:��2�f{�.�Be�	w�Q�jE	2RE���|�L����tI~��)PH~�C���Fr�k��C�wF��Q3�rɔ">t8�s6:l��S#<m�>�s`:X�g���z<s!G�~��>ԞƸ����>b��%-ܦ�"�#F6\M����Q�xNK���'���3b�^ِ�4O+���L�S)uR��{�f��߾����2*����n+!x7k 2��XfT� %B�ֻEGǜ2��?BM3D����su_���+3kE5)>�"�>�^�jQo䇯"�2��j��J����ME�]fa)��OL�$=%@i���O܀[�n�US�<(�O����ss���P�ʑ䈭@���d�k�s!�z6�T��rt@�N]�xAK�Z�?%o�8��P.t���8��.�Ãbm�E99�	%�։Ěҧ ~�f��� ��z��>��fg]��ڊ�����6�&M����-b�w���Ϛ�ৗ�ܰ<��Pe8̰Нuu��_�l=�0@�X�zQ���?�_U�������xV˔Z_�ԷZ���|����bh��
�u/;=�1��1i�d�oEG�Gq��وDP��1�s�*�A��b4 �[O��KC�bU@��C�r���J�����,=3.*C�;ѩ�F?�YV=������b4> �d�+�l<�8W=��&)��L��T��m��_���Ǧ�tl���3M��Ʈ�4���r���N�Z�6U`����TkscQHH�M���J/�j�'�C�Gs�|����9tς8/h�Xl�8-n��^�HA$J;�B�.so7�&p��"\���S?5�R��Yk�n�
�Y��TF�S�%����9Q3�t����>O��I�}��z8~�PG�u�O�4��x}O�&���?��$�Ԗ�+�Sw��\
�I��#�E^*'�u?�*��'#S����[�#��I�^x��1��]Z�o���g���5��~! `$���Y��a�X���F����Os'����^0s/I޴ALʼX`^�r�7��~����C�'q ��������C�hf�
K��B�Y���WkiZ�Qkk�Em��̩F�Wmb���g�	�ϣF[��,u8*�r�y��W�Kf�)<���lX��뵗����.Q4v��$~lƐ���<+ �kjT��b_\*�ï�F��%4��^<,���ri��Wޤ`�!���CYH��m��T
}�(���(�x[���,�-y0ax��ޮ�<Uh�H�pͳ�#��5��8YQ�H�=�8�r
�Ui���NВ�V�+��vCed����:�MhdE����b&ך��c=ru��S��������f��	"-Z��cB�ң���s+:��_�4d�t��'����"(_��*���c)4kя��m{h*�_���3]ݍW	�
4�7h¦hK	Oe�\j�V����D����e2�PJ�ʐ��b��TV�/�R�,�TS�+�]�ӑ�ם�D9ԧ
���)�Oň'⢪	���C�6�/��ɓ^]�Ma�.7d�6��۵����m��m�����O��d��TR���� 8��o԰r��k|�l��`�)��T�a��d��&%�G�%ȉd���u.M��gx�������ԏ�W���v����q���ü��$ �Z=�0�D�����[cx�\��y���U��h~5�?@��c�Ȋ�Fw��{��Us��g�X��s�w�i?u��/�q�-�%H~����پÃ8%��J��佟��V����	�>��:����`�M�N%���S�'��@��#��_>��o��X�}�X�n�&LRpK�B�ǯ
�(3���x�وje���z?�Ң��<{�g��z㙆\��������0H���w��^S��Ϫ<������e� .�����.f*R	���Y4�������c�;?Ғ
� �H�➨"��4�w1��
����3��Jghڗ�R�K��f�P��|��K`usF�υʭ��1�}Ø�����p��Z�<AD�Ǖ�Pp��a��Ԭ�V ��p�O�1p����|xv�:�V��c��4ØP���\i� z�������?@�ވݤ.ɶ;�n��V�g�<v�Kެx�i%,�9���M��z�Ӟ�m� ���b�8����qK�`H����O��[,��&�r����+g�Bk)|L2��A�� ��-�Bh��u��\��2?
L����B\�w3�z�/ +Ɵ�L7�f���g�Z���n����i��C_�ߩz�
n_ˤ}E�i����(
�~����:w��1���u����"��s��,�W��VA��@���	�z"HV:�a��Ɵ�vg�j �i��y��}�ZY��Ӏ[� �ǹ�H�ܐ���o׉'���To|U�?*}A<�҄2���1+U��⺮�N+���-|p�UEJc��$!w�yx_(a>�'��4-�+AMMl�t�'
j͢�|a4��jW�u�Mh�_`V�D6�gm.��!(�Z�̀���G�3�T+A��+닽�J9�ի��V<�'l�aB̀(R���	M�M��eW��A:����*�,��.%�ǂ:@�]P����t1^#E&t� uâ������f�\��M16׃3���'�:[��� �O��_B�5�)�����'i�CZ. ˿�cR��u=��p�-��^�
���Y) JG3��CQ�b�6�'�&+`�8b�*:e�ں����3��Ccm�s�.���A�E�(��@�p��糫���L��{�LHj��IZ��ι1�2g}'/�Ms�x�q�n����˲�<�8e�YW.��`�SQ�ȱ�&Kf�ĉ�ؼ_h��/_:�����[�Dm㒄����⃺ľ0�=���[��p^x�> �=:�j#-�1���H�j�oBG��/��� �	�M5	��6Uk���z_�����H�
�GT[!&Y����OŋM�s����1�Ĳ�}�Dj%CF���[~H<�y�U��>��T ��N�M�n�'�w50�a'���b���8��.Y��f$9�(N�F?�6��j
�6��ػ/|��5�����B����:i���|J�+�{؞�f� 3�G�RZ
�SW�tT�:vsC`�s�g��
�h�p��a�`sLa0k2b�uzP��N֝b���)`lg�zcQ�E�Z_��?S��
���M|���	�Ӱ�ee�����)zx�W�
T{o���E��W�.��v�>{2��ds�WA�_>�����k#}0�癣�Ԅ]s'K�c�s?��m!=��'��N<ާ�Q�����IEB��/�HV&ƦH���d���Rjx��-ýg�}D��������8�]9�)��u`w6MX1��j9M:��h�8I���qh��?\��r����Y+&n
�J~T��h���7J���~C#&LX�AB��\g�TTY�-��:XF9�j���.{h4�}E����ô e1�=�ύp**Y��ǵ���cH�J4.�0��c/�Y�mt]SK!ř�]]�0}�r;$k5gO9�o�Է/����e�@~t�Jݩ��F��mZ���z[?��j.��?)R+��}|�����q܇�$��k��_q"����@h�ҤU��-��4�ȯ�2(ZՔr/ߛB�=�^�SYE-�iR}C|U��=V�Ch��*��q\]�R�t(,T���5v͓�,?�e\��/��1���}wӝ��ƫ{)�)���Fd}22�^���|����bȔ+,��k�
��s�g�X~(ǵ<j�.z2�,�aEm�~��L?I��]3Ex��;����Ͼ;��!NL6��m�^37)7�	���������{ݴ��Jd����k6���^��%h�g��d��$��զ�W�����PF���/�R1Ec�t�#��73�qZi*4S1.��,��t�̝:\���� 4	FE"5�O��U�PD�oϋ�v�e5�À�5#�=�8u~q^n)E�il�W�d�Z��os�O.�U�c
�Ԥ2���[��"3$@��Jz#�A�s����o���WSnirArg�{�ʌK?��{Խ�����Tw�RX�p5?�ų�����&��Jf��K�{7l�%ngzy���c���3�ã�_�~?\�R��r���@��[=�[ ����n����@h.K����MѦ��Bsޮ������� ���;0Q�J��0-�,Յ�N�u���l� W�Ҧ�U��߬�1�*���i�W'�JM_�k�� {O��S�n��n
)���Ǆ�{�c�#b�ߎ�d)��>K-���J�U���p
Q�m.��gn����<��`c�$�2�"իn��,3�m,���d/�����^��JC}�Po�$摫P��0�ݮwkԠ��+c�?4����(�`*�D��޶zGA���T}�ȹ��7���-,r������!�z���ev�?��_�tCfʱ�{#����)�\�ʚ"��|4�d�A
<�stp�V�,3���עc��w��/`��
��,04Te�Ua��t8��奜j(�^�!>����SyP����<�j�w����p�u�=�q07~�;󓅣Ħ��ir{��c�Yk	@�|,�1���fUu�C�7i
���L��
�H�h�-��xdi��Z��
$�wW��S
�/9���Zw!��QJ�Xf�=�y�8mzA�}�F|VA`��~
�YНȮ`�O���G���(Q5��e���-k~�9�,����V�;Su��3J����3k�O籬6�\������������'|u����i�{؊¿�G~ &�X��;�r��`#9�����~���h����P���	�m�*�����8vs +���PMP~b�Yћ#�e��m�֣�����)Bw1 mgֲϯ\ L\?k�s^��݋Q�K�K��/��Y�ch�)x���~Z
nz���6��Tv+q�8;�B4�s�&P��/P���a�&����A0*
]���O��=$9[d�� )y]��$��^ib��g�YXU�㹝��[�y��m=w���\x�
��Qiu*3�,�%0�iu�{����E���z�g[?-Ƌ��e��{3|AzKK��j��u�%�w�5U�q�R' {��IXg��
�1�!Р|?1���r#���EE�qɭXS3�q�(�{��V�'��PoY�<�w���-A�p�A O�%��c�Ե�F_1��Ef�����[�Jg;$z�
�������Ӕ��m^ p�NSȠ>�Re�[�Hd�?_BLov'�s�ep�+�*�y������ƾ%��d����w�!4�gZCÈfw�Y
�Qi�}�F�A�d����i5F��0�PW�BN-hI�W�~�H��qm����x�Lva�tK�:kq6�@�H;����K��b�u��O����v��t��(K!�L"��t��6"�6�x�L�'���Z�ev56f�?Öc�L��)iZ��t������pFX��3[oD�N��s���~}!�E���ԍ�uq2[�6��o��(�$�� ��_���f��<��C�M�4j���P�ы���7�;�%���ｅ����r]5S�|�pI|�)�@�����_vՈ})V��_��^���xr5�S�<��uM�Bu����X�}!���;KE�:����ӧ��L?0�m4'#����"6��`p��7bFR���3�//ʔ�z���Re$ߓBH��U���40'�	ӔN��o������?������C+�ϥ����a�Rot�����s��{�����=���� 5�?D�B"�L5a��w�zocP�w�"�Ŗӛ\nV���79n�t/�u����S�RRқ��Tz9�����%�溬>J�i���;�R�cMN3�\ci^Y8~����F�L��}�X�Y�Ŋ�F���h^(M�?UJ<'��#�Ǹ�zmE�>A<����9G���B�N)J�L�v]�Z� F�-='�$�T��#�ǁ +t��h�����'�'������d��˲�{�ל�t�g�n��ޡ,�"����؇Ky����d��@���H����gU�5�����:���Co��1Y+���h�G1 F}3�KOQ�O�D��;�@k'y��0��7�#��^��~��%ibW���&t��3�x�J��	A˪z�oKwa���@��5*Z��,�c����No)6K(U/8�6Z��#FAô�I�$�Eh�_���M�~<3�G�0e^�{�3�)�;��R��G(%V~�i������*+W4�`%���Su))�� OH`��&v��d��E��U\6�}�Q�+���q��.����{�<��3�YD��%JR�Դ��ɱU6���4�c;lY�� W��Et�Z3��3���9S�Rg�'�:�Xd�e���zt�%�m�Q����DJ5*��������jc�bfs��<l�G�~�H bI�ʣ
�蒹s� |i�Gɚ��l��n�2��T���at��p)Z�9�:�.��z����4�<�3�b�n�����Ӷ-ýV<��|>;�w������X�����,��Y"7f*Rv�F(���FrV([Ϥp7V�Z&��㽩yj��'�Rɛ�ب5:�]��5k���	HR���e|@9|ߠtv��i!/�Z��0�Eq�^�8�m`ے+Hh\�*[3 �d��#��_�΄o#��߄�4t��nYOl	���%��o�f3~$5l�T�W��1�$�LĘ
!=@�D�'��D�ޠ����,�W��9��\�ߙ㹵u�ǰm��^^�)s�hcW�����P�a�h�纒:����̤x�{O=����gj��������D��xq���F�~kWR�J7J�9q��jm���;�Z�펯����W�6�S�^�[����2�������1BpM��A{S�����E�b4�H���t���8��'u�p�D`\e@d�!�z��a��|����d;�Y��]�Z�ץ.m,!>,9X�eS� �s�`:W{y�n@�!�b�ö,b����P�� 	8W�����C+Y����w�b儞�-K�y^���9������3�?�WN��TB�4���M:ԥj�AOu�YS�Qt&�#�Ѝ�^2]�����:��5m�]oa�zH#5�]���T �M~�xm����!�9�^���JXА8ԟ'����P| [%��!D�}=3�c�P��+ 6֋U���Q�G�(QǸ����p����?�SR�xybq`�#0f�z�z�8p�{$�o�:�����abJ��k��:���s�ˏ��"#�Q.�X5[�w�j����:�{�¯:) i�'�w4:�7��J�����_O�,�8���ϐx�p�+sw�t �;g���K�j��d��w)Sڳ���Q�Mɲ.fS��d�n���]�'xW͙l!�!˭s�^�be���C���F� ��)1��z�t��
*���w�xd��>��2�`����Q�[�����e�B�ٚ��2��R���L��z�N���,�?��m	�xn'��Y���<a�yެ���M&%G�<J�fX�s�9���-��������d��FVP�#�w`�]�8���D�@�(�hsx���F��#�����T���W���#Y�#���j��݀��;��نV�#��/�/~|����U�x��I����k�Z��;SL{��&̸1�T����C���k�kW�n��wĊ���;KP���N�N�Ϭz��P������1�c�U�f���e�C�*�a�N�Ä��{��M�lŏӆ��U
b�9�uT�;���*j�m��5���tğj�>�����do�[g:풚�Y�����8���p?<y�M���V�	Q�)�:e�U�o����~�>��e�=�5����� k�&� �$��)Ƀع�h�=�n� KN[>�t�����N�]�g7U��n�1br��gӠ�b�:�7�5)ۏ=�Z��)iW�o��^��x�"��Y���#7�;�LLtG"0�#�!�|��K!t�=^������U�o�5?hf�5�?�)���sJ�K秬QsNG:�[�0�l�(����֤����f�4׽����&t ��KmԺ���i�f-��N���G��RmY��?>`�og=}�?��f�Ӭm;��k�wm���!����{Kf2�'F�tF ��[{�j��r�|F!�W��İ��}���W����Ab��G��_��)�gq2yJ�a���hF[+`5��"��d���7ͳ9����1���8��-<>1�<R����EQ�>�,�����&L�u�ެU?,h�t� _ưI��\���l�uG]�w�?�2���m��y�b?f'-�;�&�Y��S���H���u-S��ͯ�������
��������ؒƶ���&]�($��n�~;���q�/����p��<�����'�2���|Z_�͟�0ףJ�{5��@{;�iK0��LF�-��qe�C�	��X�kΕ�U�`~�p�~�K#=�,����̫Sr�'jCJ��Ŝ"�8J�c�!p�'��w�����V%Rt��T��s�X�bTc;�N>k=�Β邉�ϯ��Ŭ�..0��c�%�)��s	�_�V�å��7Ƣ����~�Ӱ�\Px@�t�Q������+߲u�a^�N%=�dՠc7bnB���(?A�z��	�'']q-6��ϡ>)���'����N�*c|�z3J8:d�ޏ`~$!h��w����6V�J�\y�
,�i�`��a	�������h���؉��
,J�c�蜊-9�.{�I(�߱��ȐH=�ё�gx�|#�{H{�a����s9<��"���*���ɰV�SǼ3�g6��ΰ�/�w:0��.돴m^���7��<2�doG�p�'e��G#�;￪���t���0��K�Nd����w{]�B��|��F�wKD�.p��Y酵tX5u*�k5���R�n�]?d���r�E�Ku"��@�`FM�I�ꢸ#����p.aN�3��N���������᬴7Gƃ7Z{t��F�t%-I��q�X�6?@�Jn�yR��@p�@�OƙX����L�ܜ���1���K��G�Vt_�P�N��Ai�V��;��:��v��ۨ�7`�~p۔L���	���S-<�-*��#�2��-�aC�4��`�t)S��?�S���O�N��`MG�����|�zL=��'��40ZY0�z�F����0�ɧ��h�j7y���Z`r����VŻ�2|�%�D\C��<s��i(��U�eVV�L�׌���軓0y�åWu�Mz�ޔ���<������D'��Z�@Bk�Ƨ�<F1�`��;-�[i���A��v��֋AB@-�s}+=�,��W����#�����l���5���3'��ۋ��k����Z1g����R����fO#7� Y��!^���צ���<�W'w����>�x��W[�4cVz��2'����8�����z�3�b��J���;���3��n]3ջM��Y�{�x�t��w׹�W�3��#��t^WL{4�j�L��U1�)���/o��o�j��}^���å������e���`6-��ݵq7�DGv�;*uG�(x�'�NΗ3%y�e{�)���� ��H��(�O�ޠ�:��t�[�7�c|�@j]X+����X��3z���M�����L{AYs�� ���5Ͳވ�9�I�w|)�Q�pt�e�5�#,��S�"�����e%��!�'�aϪ���6�+�:�e��ȹBB˽��gt.+�q!9�B�q��4������ ~��>���2��	t��u����v�zQ%i�m�4ji$7~�9=���5cHNG|5]��n��i8ظ�~��Fܶu���L������paİV� ��g݃KJ��?L����w��O���Ӊ��m{�T�Dyh�J��&�6�x�6�L�-���$�����j)�h��ԚY�v���1�p=��~flIF����0~�)����,�!� ���w��LB'i�e+WW�)x��#o�N�MR���\��ˮ(�,�jם2ƺaԸ���+W<㸘ܼE6�l��n(���/-B�Y_y��m��H�Me�`�B�P� �|DCdj��_oj�F�y�_�?ڭ�=\��^6ɹ�V��ps��ߙ��G�7ĕ[ji+%��F�m/�.�Ǚ��A�I�������w�>j"_6�y��|Co�4����ޡSNi�l��u��ɑ�Vd<^��Չ}�7�B�Q׻�t��閨�{�k����'�Gbj�3�U�z��@�^%A���ʹ��=�o���T��u��|��&"^B�D9�r�G`��׶���ȍE&��M�Z�����y�fC
�G�����������GY�x�/����/�|>�"��8�����ۧ4��h������UW`h,��~�kHT�����E?n����@"R��;���F�����#���;8l���9(���E��c:��,ϯA�H���7?΄�s��ik��:�	b�T�?�:+���X#�O�h?�#��S�?(��S]lR��#��U
l)���t_F�8;��-����V\퓉cVA'�3nx�2�YڻU$RN�.�y���1�w�����o�s^<�q�h����7\N�a>T�2���g@��_\��D{��pl�J���ی��2Dc�^����h����d&�.95�-��\&�nBPƗk��l9�#�8�{\�a9�P"M�*��rh;'���F�[?%���{n?4�����O�8:�S�cM.s�f:j2P�ɍ�`��XX#������_i�����IC
Hi���iRW������pD�kd�qr����<��b���uʯ}��^�p��#m�l��3+?��Z�uY��a4;�� �>/�y�Kl����9u���H�Q��\r��8��}������_�C����f�:9�jJdE�S����v}{-/�+\}�^� ����\3k�8�x�L(F�~���8�F�8�}=1��)�����.�^O,�{S�:>�t�D9�l'ᙀ*�_9m�m��'�ue�Y3Jl��/�R��*�N�$l��å��!�,�*���c�
�%R��F��a�娾!E}C�7���-C6K+_Q	�me9L@��޽��1�y��0-f-?�����h�;��I���X��(w�/�N���[�w�V鍭XD���@3�l��D�c�)ok^̓ZZ+�R�o,�1�j�3M�-[;B:��4���Ү������s]ҷ �g�UT��
�Ź�����c����E����2z�~��K���Rk����|Oc*Чsi��B�,��4���ucM,��$��d@:{h���R��<dF��M���ڍ.��ϟ���ĊC倕X�nӿ��W	��,�^3}ű���@T:ڦ��-��y(J�f��(��r�o��Ϛ]��h�̧�*�5���S���W=��&¬�!z��n6�b��l�Z�hA��%
����kZ�����Ȕ��򯇆�����Bvڽ��6���A�3��l��33��*0�]����1�=��+�<����]/�k7ǩ�`��jq?L=��N
{�hJ̈́i��	Z94hÛ�Ie_&�bj�S������o^������>7<��@�\�B|���Rn;�Y&�eꎖ�B�l�����C٦�����g��ó�QE찅qҹI���\%�=E�PZ1M�6F�m�I�ei���膩pȅ���JH&��LY��yQ���D�E�t���n�	�K���X���%��3�<��
k��Ty����Z�%������ ie��>�}����0Ϙk�/|'z�;� (��rs���kx��;`�&��~R^�~j�'���Cd���K՝�����	G��_�h]�P{1�j�`EI�n��8,a�v3e�,��������-�
`}��%�	��]�F��L���!���(����hQ�џ��-�7S���b��Z�:�P�ǐث�t0:шa5<@�Ga㳦L�b�GgX5Kܿ�����ҩ ��bڗ[7N4 �����!w��U�l�ó�Ӊ@j��a�go�,ָ�t��W\�������8pz����wlC��F��l.ʅ���(���������0F��b~�3(n�N����w��5�.�O��Z�:ъ�A��-+NaS�����Oa\|}�锪�1�����(��g���h���8�D׬z֛$�F�?\�G&��k����l���\	9���5��%�J�{�}��n�`b 01�I�]���I��}��Ro�p)W�ʩ�� ў�L�mˉ%���'Uρ����n��jʉ���fs�L�)��Ys) �}d��`���Ֆ����p��7`���ӱ��Os[�Ŀ�?T�19s@l�+�9x��m�j�ԭp/I�W�
'̜II�g��1n]��l'�&?�;�΍��>T�@B.���)�3�x�7�c#�W�G��ƴ
W_ǧt'#���]�Qɔ����A+۱ڢ�9�S�ݫ9���U^qޒ�ڨW�*�ok���ҧ{s<�����ƭѭ������}f%3R�6�Z��8��ɭh�`41�ga���{�}�۫��׶
n0�q=�>�WS��m����<��t�~+���H��r\g=M F3�<;�����S{��*���h���,j}-��X�G��NPg+����	 �?Wry��X�4V�{'N�>��8�o�@�����9u���L0[�mkٌhQT;�"�Ct�QAi�9(�--�-����.�Vݨ�j2��(���MR�G�{�9m�"�II����������-�8�V�M�$j:˥���@!;�9p�М��k�(��w����-����
�a@&�Y����X�j7���<��H��,>c��������W2#U���-n+���ְ�;pV�)�AT�2
=���*(��x��?���ֻ��O��;Mາ�#> �J.r����7������^U�;Ԭ���BKIR�r��)��(	2�&{��Z���ל�J�M�k�7���i���C�)�K|t��I��/G91�X[GF*���7ڒ�1�M��H�@s�# �؀�{�|8������֫�[��ڥ�����3Z%o��ӧ������ǅ��w��ڏ7�{���e�#�YCV���'ʎ?��y$�h�����R8⁹�WpT�OSe]h��S�D��csx	u�gն��HE�Y�F]P��@H����Q��9pSd<��^�7�^�u
OUX���G�*+��N�����Q�No~:{�u��	-+����C�F��X5�e�,�P:$T�M�f�mh[$�{����
�~���X�;�=U�%�~}nj0b��X�>���[�4W�JUt���	��+�a�Vv%M+vת�D���[))53zYv�9�֨ �ݟg:lB�#�?9{�����S���K5=���뵊W��⡉����i��i�p���q���h�U-�{6�_����k��Wz�V��yZc��	�L����3�`l?|����ܤ��;�1v��鑝�u.ۚ�����\��B���a@V1��x	!�*F�L^4�A������Y�g�=)=�YJ �˗W}+�=�Zc����MmTC|3���G�NGjw�[5��M�b2�#��]�d�0��
���/�ߞ\p��>��[�%�w?�@�5xk~��U͕��l�g�b'���1��TQ�/X���V��&�E��9���U�ou��z�>�$�m���=���7��wm����t3�=�F.+ߎ��^��-�]�Qs�����'RxdJD �����9r|�쩡:�}�]!���a�lN(�!~$Vc�WR��ࡥQ��h�p�.� :��} t �!8]��[8hYɢ�#q��<���)���=�:/�`2���lʡ����lzм3P�Cx6V�� ����*��uK'���dU�6���iL]�T㑹hے�ے���?��;��=�7�E��`��HQz��RU�I7R�ҥwB�*��"5�&E"��@(�R�& ]J���&���w�=�q�';;3�2�]wY����b����p��������ikHh����Ms_Z�dxz٠+��A��@	��E%Z4	���V���ރ�7o�-��T7�d�o�ε���1ߞ��`�~� ��X��u`��(@@��@F�^r��^q8�(=5��n��E�hŬ���jbp�,K������Ί�ڔ�x�Lّy��$I���.�O?#WreV>�S����^�e�_P,Ӧ��ybn�1����9�X=Z�`S��^xv�N��dOq~�i�J�������D��:��E���;��	"fq�%_iR�X&T���Z��[�k�������DΩus�h�T-)(2�v'�L?lS1(<�/�^�y{���T��m�L?���e��>�)Q�w��Tc�I�"���o�Ϗ�X�&Z:S��-�d�,�&�.�����i��Sڠh�8c9�����@�j���,n�&����Y��F�_�E&��?^J;���}�aܩ0`0�����F �{(0(�D�ޘ���3iO	-c�OSS7���q��7���EMXA�)��FJ�ݨ�Z4�T��r³��Kk�mͣ���0�c��g�k��l��P��U[�	���?�"\H���Lp��|����o[��9���P����#��H��a��s}���m���F3V��<aۣ�2\��(Lz�+\?l�� ֚;w6��� Q�?o�S0�pF��J��k\�Yf�K~��T-�ջ���1û]�_���6ߛ��<���:Z�o��������j���N����z�������d��n�J���B[�(��_(��hI��A��z
��6>�8�)��6�2)R��(��e��Z�=���1f���Ğ�l_)���Y�1����v����M�8�����t�n�J��3�`�2��-]�Rж��U&Ƞ�5�yG9��v畝^GW�[�*�f^��������?����$�(S@��x�7����>PA�6N���wv��,�}�J�,�(!nB����@��]5�Pe��×�]���1�N� D%,�t��9���6�6�e}���u���N������(��ɨ/w7��E8|l3҄�˼���HNUc��/��ߏ��!$��k,������5u�Iq���"�2�F�(�D��c-7Kk����9	�����,�N������<'eNH�Rf�ը��?��xq���QEc��%��`�Z℩�}�?�9��Br�l7��=`%�}K��^�7�]���#⧩.������"�m[��O��3ox�s��}
R�@�J�D�C��	��*���#�Ԋ�à8/��`��f��������R��W�^8�o����x�g� ����ի��Rl8M,]W����f>���΢����k��)���@'�� �U,���>d��A��,�Y���
�+;�,����<���%����g�cT���8ͣ�/��d[�c��XR��_��k䪑��T�/�1�/լ6XՐ~3�E7�¢�����ru͓ϡ:[Z�%� ���	�SWp*:��C-�펵��j��ů��S³�MY�0�v���'�Tp0/ kJfw{�c Z��� �v��)���h�To�����*?A���4����5�M�EEw�o"�풵���T��,[2�.e�nJ9F��p���&��-��)�jPI����|�)��|�e-��'������hx�ّ�!"ɽ�O��G�C�mOuGѽ�$�i��*��)�Z���v���9)��}�Ȁ�1D�/{�4�17IU�2ń呰{}ǥ�#���)!5�k�� ��c_��yF`�[��?�����SQĪ�����r�)�}$C@Mxn�:�^i��U8<�������oE��ڪ��B8 ����/0��7PR]��h�j�Z
&j��|HN1f��������ס�k~�JIۨ�
�
��¾HA�L_p�rG�����S6<1���X�_�O���cI/��Z�r����V��G,V�Z���m�r�vFvl2�'�<ܜ<��o��P�%T��#a�lrv�M@o��R9%���O@?�����Y��}G|�Ai|I�����I��d��+v��Ɉ�a���V̰�/�����;z���A�{Ӡ��w�4����1��-$��A�ʭ�0��l�^�W��~�8+�`���n�4dZ���9ʠ��o����9H��G��J.��@���ז��5�Q��)���n�o�3�.l��I�"�YX��z�D�q}�2��ֶ�&2D���_��D��E6��q�[��z��N�fR�.�n��nܑ��,h@�A��Հ�t3o�ɲ�����;�.��Z�'
�,�=󉽈�I�y�]}�z����(���{kM���m�ֹ��'�у��ͩʫ�{�ȽO��\i���Ç)�r��v�V(��A�颿�m���������f�v��Oߴ?��t�]�,�_�ֈ�o2�;�Q�c�������6�z'Y ���[�*�r��olB��{�t��B���8��N�ί��+�9��<ۣu^2�#]���{G[��!�: 4%B}靍�G��z^��d�>p�����@�3�\p�7s�v���xz������ͦCzC�����=�XZϴ/"|[�dF�v,�t���عF_�_��L��n�if��5�2ު��C6����s�ħgQm�nm��)$�e�t��g��A���у���^�$Q�"��;C�ۍ�{M-�w��_�=��4�,ul {�8r��5�?
���{Ԓ��͍�;?C8"�>Ÿ����R��꿯K,}�<4!SDV�`�#�:4vIc%�O�
Q,s;&d雭��SL�Xi�ö���8vF�6g�=���I@��l+���/���T����4�'��.�� \�	If	�|6ç�Ȏ�F����XG�`���/�Z15�0{�:��UX�[�e?r�JewZ���@���3�_��2<�n�S{��m6�Af�	E����ߥ�^�C;c|tRT/鴟�q>���P�q��t�Z��z�XL��c�غe�vɣ�RZc�f᜛�)d2�p�Q׏� W�B���5K|��#�L���F*������|kKj��N!���n�&=�`��X��oF��v,,�����mN�/�Q��dH&����B����=|T�.)�9Bf���S�0U]	(H!�v73�E�߭9�G�_k�Z���X�0lU��
�L��}�K����6_���E���6�~D�c�ye�tf���p�P���+n��Wj
߶�к'ac��qλPC��� �?��,�S�X ��Ai'��C>Vu�8�K��z/�%��8𵫅�nw�EW�3��f�9�IP�$���Go�/�m{o�����F}�g0�)�k�c�åLEP��GW4�;ry�D+S�
��7e��8_��b�Ry����4{�_k_��{�B
����z���J�l0�]���-|/��x~?A�;�^��~�(	�F�z���G62�rͦ��;��g̭���VN��/��h�o&�d�^��.rz�eo���g٤sM�C�2ή+Y��[J���t(��=�)y���*w�PݮIMQ������j�������
Z����$�dLL|�[��*0�I��C�/��Yܚx_R��kv���}��h�A['�F������0���h������Z+���������4�޹�P��t�:d�:d)׭�r�c����{r��X�E`���85�gdI�����W�p�p|��ʹx����@*���,R��;jb��ZdL��Y��޴C��a�;�B��
�I�	�TO���>��ߩ���bY���mZ=��	~�PdˇX���4s�ڼ�w��{��X��f1���һ9o�3��K�岨U�
��T�� w��Qv�dg�.'59w������������:n��y�jA|<�fg�)o��W�ʙ�.7�*�j�.j*&|d�w���Yb�R��tF�s�o��Ů[3"��Cv�_}����3�X	a}�C�]��� Ï�+��(�|�����{#i��]����g�.7��i��^i�	�@Jiwf��O����n&n��L�]��hn�
�z�`��#>����k�ciI�	:��-��9�(|3}'�����W`�~m��_����� �� DS�5ڣ�;�ö�(뽅��׋��}�vYHv`��n�
Pu�[�Yr
�g%FF�T�{O�����@�+�������R7ǁ(���_�C3p��>T��t�P۞�إ��Gc.�I����l,��a�z�"��A�R�Oضv�|{��B&J`���O��K��KN�������8�� �t�q���\���U��K�Y�AF�?�js[=��-}���Ne.T�?�q�i7��xEZv*͒7	�'A29�c�:m�#�#�)�vlշ����ii�&c���"��M2��@� i�,�3�T˯���*3^�wJ�ė�[XT����'G�M��C_��wk����%u�{_�mP�r-i�!`l�k�|�s� �HK�  H�o����������u��w-�ӬE�3ya׆�z��^&��,��U���6�©�"�m�/�Z���L�nSE&���~�ʏ�g/0���)�-0�s����Uʶ�އ��aTf�ȋ�9 ��J�A�ݸ�%d�Rt��S�"n.M�a_�R��B�i��(�GG�~����n.�Y���YmZB0�@�����О7�a2�Oȕ�ّ̅��Q$�+���%�8�6a��|\�X��^��K�hՌ�s����8dI�F�>�DmW�d����^7o�41.1nf�v�TJZ���>��Mf�H�I�Y�@�|2N7Zp�I� 
_�>�2�a�d}�!_/�B��:]�<��վ�W2B��.I�{�
���9X~��j��AWF}c���uw��p��1�Db���9���eb9}a�6���l�<�j'!'#W� �l�U'��A?Ԇ�>L���P�|k�~��b/&���I���g�lZ�-��yw�:���`�T������{a���K��g�'���o�uMCa��\��i��C 
����x�J����a��wȍ��i���.�;��	בi?��
������_qњF��m���^�\Np��ثu����D߷}�-22�K��	�*���'����ђ�4XVw/Ŝ"r�[����Y�tu+�W��|��o%���ӱS���j��(��X�Eu��1!���m�W��Af�f7��,���&�[oz�W��L�o��g���+ߠH�R��/����䅰o_�s�����0�q�V1-����s竿��z�p �[�3D퐥G!���k�P�v��n>k�����1Q�.��QCԖ�a�Z�#��~U�R)���Iz�F'=�/{C-)����}'���:�m�؂d�f���&
A�l�G�u��i�M��U"8^�y��N����Md%C�g �G�
��E�V����*�Dt�H(��ɞP	�l�Z��K�4��x	]92����))H�3�W��*g竽�=�dO�������V�,�م��3z�;��$8"y��_v�v��%��cv �gsr`���/�sk�"����E�����i��Wv�A��Ӟ<_�#��_D�mӵ�oǣZs$9�9�qcW��OZy���~wiae���D�4��MLҍ��Ѧf����3b�&�oj�^j��kt}U�ؖ�3�ݦ�Q˷�)��P�NN�g\�����oTE3��%��d3M������tᙓq���|�����gY��%�Q���N�����q���j,�H���us���,�	�4����k���3
T�p�����/@�)�i�V��4L����0�ȱ���4��ɹ�7Ebvsz��J^R���/���IHp&Sy��"�f�Uj,�T$_��1�P���X*����#dBl�	�]ʬ�אez�3���_��(I!��YT9�
� 	�V������ ,0籖I�q�\0QF�E���H�q(e�u���9�8��_I�N����H����SE6m#����?{߳W7{e*��V��tk��R6���<�ow!<�,�8��L���[6�Z⇆�OH� c�n�L��[�CZ�w�Y�Z�2�%T9?�h�෬�3�od�������Q��T�^�p��:���������t0 `�j�fCtA�x��Ĳ27�f�%ɠ�n$�c�����;��0� �@qo�#~]��0��
�G9r���:���	�;��~�b
'Y{r)	=ӫ1Ş�]����k���X���^kw��� kn���$�$������k&�2K��.��	�@�U�=2h&
��Tϕ�nf�u��Rc%;�^[��Hz����F�����VWKi�%�y@�DrH�?��LP�4u2k�^��������a�r�\�����~�K�dF��)�%���e�떯f���tZOi��U�>�
�Ua��\暈�Q��@�ݧ��L�ZE���yaSн[CS��]2���a�O�B�e`7=���=Ɣ}ՙ��".� �v�U�KF�ս�W���&R��,���%_�U��6:���'e\��*l��]�7�����@m��7{S�k��c�y�o.�N��/4a��&@�4뷃�9��Ӻ�V؏V��K�{���5qY|Ҕ8{�Z]+3Lr�7L�"3���������-Kꗖ �/sa":ÈA�՞�(�8�xگ�oD�$���z#v{{Sba��:P�a�@p��#�v̆�E�l��y��6h�-�oQ�08*N?���d픉�b�"!����3\Mɫ1R����x��D��8�q���w����o����k�/�Ю�55��֧RϾ��`�������Iʖ�lHgf��}�5ϝcs
��ۣd#�
%A��hisgj��󫘔�ڳ��ƒK���ʓ��@f�nm43��\X��γ�w�Q@�j^|�+�u��5$&;�!�1/�b[���y�]bE��~���w�O5
�D9B�i�����f 1����/KJZ���w.,�(�	?��J�����Jb!yv'���;Å�(���Ψqѻ&�>�W��ʍ��YEEl�2��i��;O��S$���gR����b/�~6�S>�}&|o�%���� �_%a\I6�N��&I����O�U��A%�w��f�W�, �wˀk�g�jy:����ԯ�	�A�`�,���Q����>%lhp�5�����~�<1�����G�B�+��r8f�.]��!�B�q���!�,���E�j?m�h���q��!T7�?jd�ճe@��;9Pe����pw/���/�b]��TLO߿Q������K�&���X�rfJ���)a�읍?/����"��,+��T��J��)��+�WH �C(���n��gpN�C��+2R+�(��M<|;��@:ئ�������y�m �zF�%�Ff ��Ϲl��h:��ì��@���_�mޏ����)��߼&�z�O����rHt�k��u3�N��V�-6�� e���ʤY]�cxJm1l]b��j���;4��UNiB��;�n���c��"�WM���f���͇Z�_��w�B5�'Y~лZ���I֓��'�O�@K���:+�&ltr}�r���%�H��Q������,���g�ł����t-$P��IP��mڐ�0���<XTΎ�>l�q��8��g^���\\<k	Z7�����R>6��hWN⊶?�p�9i�䷚Ge)�K~����4I�z��7�ow��5�k�H��Q�2U�	���-�v����"��%�����Р�tK���l�Q2≮~�F:�-4�
�$`�V�*�?ܸ��%W,���D����
�i3���i���{z�vıO,`���s��.G
��`�6�����⥫X_y�����Ԑ���d�*���}AOV�t�����4l�?J�h,�Y�č��1yk�'��q"I�ii�(�`"Q���$�R��覆��:��t�vO-��ysi2:�������+����@�fӛ^�������!�mH����/���?��x�,��ͣYg�\JV��B�D�ۃ�8d0Ŏ��@4��(K3ס�ixC�u ����o�E�l��e�h������	��)��ވ|xP��='J%�3�����k�!��K=�W�_6S�`��\��� �՗�?h4t�yk�s�.6���7�r��ހ��;ǎgN�K  @��$�z.��d%=��ҏjҸ�&�&o%y����]@0S@���)Uj�voE?d�y�;Iy;�pH[u�?��� � i����:�t�z� cW�y������Z�3���S���/���t.����.�J��t�G��*�j���Y����/�G�>-�%���1]w��]Vi	����7�p��ap�ŗ��:��x�w��ԓ9�����E��v�R��,���d:ҁ�$���O��K���5)�����?���.���Լ���@c��';.�E�;��r������P`�q"��L6��z��&��k�L�g,�ɮ��]X��u���U���b��7�݉7p�P�1�;����5��WBؾ�(���w;��}�z��Z�u=���M�eHw]�݄��[��З�κ��!k�C���y`=�P��	[�x��16mIq]���ž]D@ u_D�_j,���i�m�X�(�b�]�>���5��j��e�;t���(mj7Gy`�@�ӝ�j�۹Y{����'�����)�����''��R� �3Z*(�0���q��>
����>��9�i��!���Է�}�*���"� �I־�=��Iߏ��;��P��;��Э�.�W�!��ީx��ɮ>}�4�3X�i�~%G�a:blU��:L���|]d��9�:���d�aI�<u�\�-�����X��V*���/�o_V�a����O�Z���y���[
*��B��P>T&��߄�K�#8�f�Ї�+b���������x�����8 s�4{�c���ӱ�L�,���Z�v-�6���
i.2d���!�_��i���oG�g���>a�'�
5���� ��s0KY��K�j�����DJ�*`�^(h�4<�L�;)��h-�;���^�Iß�u�>���|�>�J,�rc�~X؍���k��x�s���m���VA�7�0��kHz�ka�<�sNm�R���C)���r���HMK�V=�
1�;��܏���#���/\_1�>&DQ��a
��]��UK�1���%�e'T�/�����k�P�Vye���MXc:?�I2���{��N�f��A?�/��'�a܉��*��&�ۋ��᥇ӌ����)&Yk�`47�G�I��X�/���dT����˵���XC��O] �ҁ������n^V3�'��)/xX�=�~ �R��ppA^ + CP+o$��C�]_u�\��^��|���%���v�~��M-6h�ɞ�詒\�ŵE)Ƭ�p�F[��F�mR;�y���K��[��E\4���F�KN�����f���ا�]~�3�Pކ_�>�PvsP�Q�I�7�H�����%���'��w�~0,�,�Q�m}�T��+J���r��B��!K�C�?߫ 3 ���bi3�gL�K�~S���c�| a޻��g`C�U��q?(�m��F�<nX�&���V%�R:��Q����� ��ݥl�S[;�k �2$�n���E�L���[�I-\|P�7�h�( S�~��~,��냄1��8~Ӌ����( �4U�R��0��EM t�|h�@������*���g��Q�1l]�e�Գz�N@FK�J83b�܍��h��x<�i�v��kW�lv�t�ܨ
m�m���{��,��E7�s��]�v�x�����]���2F���m.��#��Ғ˹����ߡ��T����U�h���V��Z=��O��yڅFiW�C�56W�>�ÿA'AI_���x�B:D���.�����l�o�dk��ꗚ�%�Ʀ
#�$H��mQ?$�	�������1�0.�R����>S���C���5�a����O#%U���i%B�Ͼ��k�ş�W_�	���K=�o�V,{?A���@����d扃��#���k��5��|F��{�=g� �0,���t�e�IB�d��G��v
��l��`�ۜO��sX����D�K3��6�~��h󩭈�����Gj��W��p,�S���1#R���
)z�d1�֠��L�M�R��2�_�\�����aj�\)S�~�o�� ��D����ڴ8$O�	6�'�8����Ɂ9 wtߝC��p@ߚ�545���������E�C4����uw�.�b���!�酪a3���Q���d�\��qt�_�J��@�9���>Bu֩"�ǖ��%DZ?�I���������)Ϛg.���.Ų\��
*�x��xwE��wt�ͅ5�O ��Q5C@��U{��%���ڸ��7��KT}��v��!�`���@6��58���3����j�T�/	;��v��4~��˲]w6������Os� �;�xT�/鏒6��6�g��N�-��9#�NŜ�]c��L��
O)�N��E�Zx�E�B6���A��Ĕ�U�)�{s�p��\1GJh�5�c+�@�
��w?�����v�z����="�� �5H� 	k����&��j�]��Z����T0�O��x8�6��������we���D}�j���f�ZӀ��O|�K.k�nc��X�mU>HOKJ�.����6�tN{�Tv��q=� C5pW���#}.�c5 �p&�k[$�c	1�w��z^$�r��P^�, �ͻׅT��O���]t/ J{�T�*2�÷�V���x�<��ޕB�3�.Di�����u��w�X���F]:�&��Dp����h��Ȧ}1ߪt�M�H�a�Q��/ܶ+�ё��N��-@pt�V���o+�����.z�1pa���CW��,�}��o��p���׍(ƏF��~�ŋT�z@]��Un��.�,z�-.�AF�Rך�;kT��5�d2�"�O [�xn"B�_�$2�zS|����Vp��,�$�k�g��/�a>i	:�ua��5E��"�ๆ4� �J��^�:���u��;g'}�+�V`�G�����|�ׇ��[�n���]��x�!%Y~�J$ӆ��v{��`�h�lyRU�(��߮�%{�úf�X?�0ٚ�7 vѣj��'��YT��B݇{�?5������+PP�*����*�Gj�_0�MPO�n�K+�ܿ?� �u9�GN8a�d���N�����S��S�������L��D{�ޅ�x2�=+�ae��B��|��:�u�=h�)/�ڟ"ώ��V����Q�$�]
��F�G�cՒ��`�"B��|��Շ�Kܜ�}%̞�G}?�T����,^�f�yʺ�KXȍ��7bW�߾iװ����Q��`��|��Nw4H��6��m�.������H��ou[PkxC]d�Y�5@`�Is���PF��A8�yO����x#����e1���q����w_srU��W($�<�JՊ�
�+�y�T��ajS~2{oV���TZ�d�_&���|EU�����T�f����U@����z���V�/�n$9�)S�J���f�c��kz�5�#]�Gȉ/;���9p����h�&�1��v�ik6��C��T����.B��E�,�;s!�1�-��6R��n�]
��w�[�N���5�ӕ�%�g�X���8?�ufv	�����_@L僡�6?j=�� w���Ir���\r��9����GJ�����m�~ׯa&���c�W19g7�}w�Vc~L�~��nA2Exܧ�7�-�5nR&A6r��2[w��w�}�S��z�yՆy\tȟ���SxG�H���=��/b����91����Q�f5��<Ey��Ne%%'&�Hݎa%>�J+�raQ~� I��JʪB���(�����x�[ŕiTUU��lc��>$����;6[�����d�2�'�'�y+�=��jzjjUm����ЯG�R:�'ܾ(��gzg��3B1�f�h)q���7��˥��Cђ2-J<�Xn��e�Sb��'V-����in{���*���j��%!Zn.������5�O��0�;�U���x�T�4`@~i'�\�E�����iJ�<�z�ڎg/[L��.<��t3�U#_��ѿ���&��;zx���e�u}~T�p�9��Hʨ�����a�C�d��%��_�'�+<
�8
���cMRj�]G��m�y)mٴ�_�ߪͨ��;���K�>��b�UȤNl�i�<`�k������X���l�Y��ҹ��`3;['�`{;���uP�L��?�9=��Q`��jH�+F��D�^M�v�yq)T'ey��[�L���u����3x�(.%���՘�����V�y/��_�^�����;m�*�{*��p�ø�yǣ ����n�4j��)O2Ne� l��9^����>'�w3V�5G?E�Vm�5l����Uv�,z�
y�r�M{O�i�h��{�����9����1{��R��6a�Ռ*���'�o�4i�$��^�v�V_'}&[�P�[�ã?+���$Ûؘ�L';�]���&I\S�%m�����b��y�	=u��Y;@;f%�!��;M�B�Vs�v����V��xV��O��;]���׿.�����g��;t�p +�'8�C�k�(o�!�)З;�z���[-�X�6Ɖ��i�rsaQ�-Q�����aˣ��_�ݸ+��˦U'+Ob��N���)t���<�ƙ x���,�4+l�]}k!\�Q}�Dq0�궧�K�P�Z�΍�1��xc�iS��v��+����xX9 -}.�j����?�� � �o�{]Z��5~��$��x`@��W��N�?��2W�%��GSF���NT0eN��w���TxݭXQܗ�S���Q�@�4V3�2�+��+�j)����W�t��h���4��8��AfE�Sވ}&X��Tbc
{{�$̽?��C�:����x����@G����2Sށ�U�Xi)}�$�����CQ7�K��-f�M[�UC��A׊J�C�S�S�m�0H���������ߟ��E�����%;Į� ��®��yuǪsjq%53a�#���&���. >�[����;�k&~�<~��8�����<��nY��n&�׉�'���N��q#�R�.杋������B�ki MY� N�V ��0fJ����6��[W{�S}}�W�X?��Y�k��z*#�< %9N��
ѯJ�CUa}�@v1s?�P�hU���� >*���ě���&^�U��~�3��r֥�ԙ��� �B/1�?j>����_.eK.���V� ���>�O�"���Ñ�U�R#��Xnϴ+zU6N�)�m��ɖ���� �N�~�;�Bd�{y٪*�+mL�է�|uB¤(�-��Y~�֞�&���g� ��Z��y���;�\�|M�����&����ԥ,�4}���q .�[�RK�:@��y@2��Z	���,]�Z������_~dj݅d�8��jߡ|��4���o�xA���C��U�-Ȯy6\@Q��R���|��aӖ��B�kݲ@3^����J��x�~d_�>�k\-^�U�^�J��o�|9U��$��w���ɔ�����[
w���}� �T;�GfM$���07M���~�E�k�B�'�]��\^��3�ϰ�uOƏ7�V/7uqܙ�ö;�[%�, ���ʟ���(�u�%m�;N�L|x!V�5��)������ֲ���u���M
�yI$�0�_u=Vm���_seک������r��`ՆU������m��i�n���tcy]��{7��l�����7���|r��QNN�؄�4\�xCM��g?V�}��1��a�O�m�;�n�iz^�u4�q�Tyh��e�t�"�=���0 �#�ڀ��N�P��+a��vG�\�~�%L�u�&�[�EF2��o��~;��)���.2����+���<�q�}�I�i�bK�L��5к7Q��%<�z��A*����4��4U��|��a��9k�NӬ�.��H�X"ŉE�(�����PZΡ� �'!�ko1/5j1�ک��YP��<��D4vyc�H��1]���bk���]cO7���;�zpПg9�M��Wo԰E8��H�e�'$D��W�����K�z)���G���j�iI��G��^b���������1w���@��;�y.C�O0�v�;���h�n�Qk�a`fs�꯭��Db/�W�"�M�?������议=�	�1�z��a�s�g�L�'7Г��G#��s��aI@��`'���/��]�]���vfƝ���1x ��P���<͵�3�B\]��u����6���s�	�rb��ۤ�������U��'#����X���s�)���>��y������ۮ��V����h \4Z��E�&	��[�Z��K����#��c̟ޞ�w����J�_O�fF�h��j�c���7w��"��]x<��jҜ��'Y5M0 �sMO%	������e����kT�AUx��o����}�$�b���N�`��co��xD���?�	��_�|j������7ޣԐ�M����b�@�?��%r�j�M����hbZ'{�\��d���O����F�OG�y���8y)�O�5?�g��z�0L3����iݹ���˝`C婙��j��_�ɫ��ټ����{��n�`=���:�����{�ࡖ�jJ��ˁͿ�v��캆�h�6��]AlU��V�Sߖv_������� �p`T���M���|-�w1кa�dd3�f����/q��7��Pe��)8
�I��OG=�Y0RQ��P���Х$��U�4sF"�.��=z��;�̈́����ۅ�30�c��?ܽݜ�5y�ձ��C���#U���	�����qm�ډb�Q{�Ȝ���w�v����RAyb#�>�6Mh���6C8|t8p-�0�d/G̞�Ɵ\�$X���h���>�~[���
�]��&،y���GU�xFT@Q
�d���p�A6	��)���_�a3ح@�;��1�>*�j��M�Q\�t$�G	ss���n��Qu{��#��?c��^3�;�Ȳ4Ҝ�,ڣMʕ�V�ݩ�����פ����nnD��o|��)<{Q%��{��e�i�i1V��c�����䕮�U��z3��]��S�ƢA��J��S��@���m�s�B�Q�f1&����J�1���Lv�֓=}ڥ5L��3�u��Wi�hR��;ZԬ_���0b]M|�����n�_�����j���D�H?�^�Q�N�m`�^^%%�����?��9/�@�5��n��5��f��Пaj���g��,��w����ש x�[����klщ4�5WdQ�E���;��( ����l1m�=��/���wf��(���x�@�o�� 1�o��NQ����G_�˭��&�8�YVp1(x�KO��.��]���	�m�S����ӿs���y~L1"�<~�~Kc�#��b��W�DH��z��$�#���ּ�cn�V��:���!�g� �:8v����Ӕ?�I-�$+ v��s%߸Π��h�KPL�#l��{�gos�[ױ��!�U�ӈ�G���)]����N �Cu �I��������nB~q���%`'������e�bq�,�&��桮��j�'A^i`���h�ub�%�.�'?!�Pg��#�I��/yacżJ'/nq��/s�
�I<�B�ȝ��[y�?/"�o�;�s%�23�O6�粒�'oH��q" ��EA�������<�����;�`j�_};p��|��a_L��)|�� ;�u���taM�mU�I$�s[��D,�03aKt���f
*B�kE���?����+���b^�/����*4I�HHšH���pSE���#�����ͅ��m�����j ~�ݎv�rEt�#���x�W�p���ߓ�!d����3-�0ET�Sj���_]�4�|`(teL�hu���4q+���K��̎����3��_���w>e|	lX1r�=];v�A���zo����b[O��?s���K#�ڞ,���`,o��}Q�H%S4Bq\�eS��	Y:�jGL$��D�c�"�x'H�ua�4�_Uk��cmg �.�a�Ɋ6��8��T
B��}�]�	�Q��	T��\�PͲ�'�"�B�f�KX	<:&��㦍9�a�9�]M����m��y��+���Ҵ0��<Y��T�M�0�K���Y��Aj�4kg��;M��7�+Y-�Y5x�>'��5�����B��P_�������b�^ƽsVM��TSn<N:@@�<�U���,̲Z,��n�{t�k��P>`�9Pq�|>'/r�W$Ϲ�F5 PԸ�C��8�Я��nF-�CrW1]UYM�q�jG���gGT�"iD�w-B� K-���gW׆�D�hE8B�̗��N�9K6�jWۀ씚�����\q��RWخ�jyD�2��O?����m�n��E�@U)<�:|w���JH�HϢ�@�X(@Pf�v4�vy�u��j�����:���W�W��+v|�3jE��>�5fPh�M�1�?_��o���9
>�;�+N���?�;��ݣ�'&����������V�4�ʓǿ�ϭ�0�m�s��>	�}/ H���G�c����[�:i��ve'/бOax�f&8��Hd�L�u�-9�qP���e���Y��2T�!9=�z����R�x�(>D_��H	̫~Q(�W�4�?k�V��Q;$0���#����v~$�X�~�u"u� �6�O�PRӥ!�2`��Zpx��T[�� ���+����a@��K��c��DL*^�]]�Z�m��!M�g9�2<S��LO3��j������_�b�hO˟Յ�J�����ޖ9��@^�T�@&��uD+���O������ �ۑcX���@����`�,�)����b�@�ؓ5hgM ���xX\���7#ʓ�K��3g@��q��)j����|�RJ�!c6�c	ةuL�ο�J1�{��؋A�Ӽ�ߋ�eIuR	�I����gT"H3#�=�!;���� G��*����_�_�/�d�����?o�5��j��J~�9�j�./��2�9���&bA�X��z"���.�{h�ۅR]r9{�_i"���}�J�۰#�����#Ӈ��	��Z�����)����+.!Ƴ8h'hw��VE �)DD��~�Q������&d���@}c44���y�!B2���Xr���Tp��z����!K�DKef�w����:.��k���*"!R
J����H�R��0���(5�*�"�1����H3��59������������Z׺ֵ��g�1��j�`g�4��$��*d_�v�+�M���S�_���&���,)���\��������5�C�Jw���v��כ�yT�U�`��{�&h�a9oP��v8<��_Y�O���@+�wӤ������숕0o��iX�he��f��M�?^�$x�"��	S�An������?��3/ѐ���G�0HȨ�
=�'�̛. ۬N#�n�j�¹�AH��q\���!th'_ǃ�K�OE�g�Q* �j���:��t�^`��]a�+�m���MD�A��l�q4V���}����������j���+��7�����46D�hA٦���U����*W耤���.���[{^�BG�Ô�$�>�1WU�Y<C�h#꣤�S��uf�4��Ƀ��6p�����2����hd�yf} �6�hy�YHR�ۏ��s4�
mH�n֤RP���6�[��,/���D�y�S�{�2�}�����2�Ě�e��D&�ȅ6rīn�yKb]N�D�D\֚�60G�cYn	&k��)�	p�ι���l��ڿZY�,�`�`jBa��חn��WR߁����&T��H�!6���@��4��]s��\��S�)4{!hS���v˾�"�����GBS�A��-��W��?%��1B�02�`Y��{v�/�5SQo~�����_Ǌ;�5�@2�G������W���ͬ�='��P	M�_uo`�W��u��4�S~�*Z'L�OMR��_:�\��3]Gl���r��O��ǌp�l�E�k�A��*���>�*��Y���\F}�t=PgC�~V�++0ph}B�o�ľ��y��?��*����3�G9���[*a�\t.ߦk��0w��@QE�}��3������a}��h%��o-#v� �e(�%���D~���M�n9�A���DO?Jt�tV��wl����O���f>���j�u�Q[�`o��	�J\[��C�?�y�ݠ�w���"�L_xS;Y��B^<h�g�s�E�)t%����Т�Y���d����W^��+��=�$� g�uɮz�鵻�go��y�Ys�&|V�\B'sx��܏MR����j�䩩'�g��K?kTR��g�7ʆ����1�?���݀�Z]�ow fzM�jwt�XfaYz/!3��̪7�z�H4��/	D��g�ӛ�#5^yʭ������}2���������,���Z'�$ѡ����Jy8S���6V�7Kr���_�_q��a8�o[T���Y�vz��ThA��o�8�B��wQV}��R���M9�s�<+6�d���ݗ����8)��[�fc���|���~s_
?�q�Nw~�T˘�&R5�F{707���m���֕lPzk�[r�N���F�C�`���6�Cޥ�S�-1O��2��B;���*ɩ�8�@x�6����@h�I��F}YL�	���{�����M֞q���ER�&/�]���Guƻ�c��U��9V"R�x�ӡ9e���-RX��=�4�lmU��G��K��T�35�8^7�q[����dO���M|�J����P/*�9Ս���v��"��y�&�f_��f<;ɉ��>��c�|j��b�<ٳ�Z��@ؾ�aW` j�t�|w��
��B��+�#��L����jsq�\ZL;_��hf�^���'�����Sh�ȱ�!lB4�������%�_�w_k[0P�A��7�L��3/;h͙M�4�p�����+�^_�����j:����]�o�Xo��e��d���z���Y��x�
��AYl��=���4�VE��7�0�-��^��Y�GUH�9Y�&��ճۨ��p"q'���M&=L�>31��!y`p��0b"�aH@W��,me}��[y��HZ:�=�C�j�;�����n��<Ͽo��:Iئ;I\Y}V-��>-Y�F�'o�{�Z@�P��1ʝ��Z�{�ٔ��>R<�]4=���@�`q�$� ������][�.��r��|��Ķ�����UDAQ�͑d�9�<M22��9�x�|�.��������~Bs���;�+4���P���
�Ƽo�i�!���{]i��V��Q��
l26�_��$�kw�9v%���ڇ�C�����TTt�ӻ)4�$��S���oWΩ�� 7��qgv�ͩӔ�)�@+S�[+ۭ��k2|�0�kӷ0M���)%�s�gM<~��n���32��/��nQ�_<z�!�5]��o�G�ƴ���%:�n�������3���=��w���#��l_4R��X�	'9�&�3,��4X�.q��cN�����R����X��О����\��h2tgܠ�i׫̈́��v��)3��8�"�z͸�{�y��'�<i	ƭU
�V�*Vj9yq��}I���	���lL��n\�S�k��0^�
���i��xP���%���@We�h�����j����Q|�x>$�N���Z�w')�
L���G����\�
�Oٙ�!|�3��`�u�X\{�h������m�� ER��kz?���~�R[��2��N|f�頄x�`�����B�ϜAn4\ʠH�t�`RЂz�"M
q����N�s?�S���}����<�dq��`��(?{����?��{+ʻ�����ؔ��ZB�7���]͞�j��~!�����w���h���w��dK�Y� *4�z�U�جT�%�Z���_���
�A����`��s�o��q����,w��W��4�9f%�Ŷ��DPx+ͨ�:�r!��#�v3������,��Y⢈Ec-TH��^���	��I<��'�gz�t��h��p���͍����;�׭��&Wʦ�3,��j��w�JTr�<���˞�!���iMm���R�����ߖ]�ﶍ~z�E����nx9�����)�S�Cr��>��ǜ�Z9���s�ZfS	N���S�P��a�zjm|*�װ^dv���9��x�9�9��/x�U�	"�ľ�&��K���&��y�T�	Gڮ��b���~��u��Y*)�ܨ�w�����K���S%ߎ^2�gsG�� ���v�Sle;ت6��M~VhY��Pr!F�ˮA�/�3h�W��hiT��I��o��$�]:�CH�v�����91~Y�K���#ô�X�_dCz�-����#�M���R�r�ގ�W{�j�9�&5����;���jR7$�#�ʞ�.|�I�j^�������ņȔ�l��mE�Mo��G}������Y�쾠��1~�
�F��O4�JyJ��[1�CĠ%�fq1�u�R-E6?{L���6TaQ¤��^�T����@B�;p�o�5��ߍ&|��{qw=�a�W��;ǔ��26J�!U�Cb�Wk҃�W�j�� G��?:�3}�Y��nJ6�yQ�BU�?F��J��Ƣ�w`�OQ��Sz)�2vfojj����}	 	fi�b�C�9�e�]t����՝��PNְ���{<��h��?���|��|}���{(���� fJz��M{k��h�[�p��i��H�r�X�Mܒ�_ ��)4>��P�S�)k+f�0Z^�)Xܼ!1�\)���|���6}Wԣ%���BQ��G^m���� ��Ge	�t�wb���/{��SԤ�%w+�/7Ɇ603Ngi�z	������//�m�����uW��.�=ϐa�����t�����b�Cb^�;��K�.�Y�ֺ��ɬ?M��"%���~7��a���c�G�s�^�G�ݝ�n������i�a������6O�]R@���Ϣ��U�i?��������[h��e{��x�c�0�+�S?���'� /���06*mą͜ـ[�! ��n��'BxFV�����fxQ�W��{
��Nxf:�����g �;�\�����[��.FӪ�RW���v�'}ʕ
�
w��;j��#%��y2Vm��	��)��lN��?g���r�u�e\����R#����ڇ�c��2��N�>r`bb��G�����0%\�]Q.��u��G[��O��v��/���k��N�ܺI<�]%�	�_���jV�霪 ~>'e��fdX{C�K�ӺjD����yx�ޤV���
���,��ܺo�����t�y���V�d�����Jy	�	!p��Z��/��^6����R�V�����2���u��qq�"���?�}[�ﯲ{�.�ȱ3i�P�g7�ؤ�� ��c�h�:Y����ˏ|�kht�;�h�UeL�#4�V�vwOd"S%/�U|{@�<^�՟]O\���M�҆=�s�Y�_��30O�J�ϩT.�վe��i�dn�
��T6���j��K��M>��yK�Ն��l|Qf�Z�j?Ea�)�=е���kR�@wS4A�v֙��0����� ��?���2�����C�m�&t��o9���N�A"	�ϼ�^��l;	ʽ�M�k�c�rU��|���$��&|̵�c@ՅI�\h�;#=��N�qU6��~�e���|;B���|�Eo-a��w=�
��
I�"�T=�X|�����D//�~í���}I����R�Q�M�g��w�mA�/�����-��4������؞�ӽ�:͞CR~��e�[ʠ*͑a��EH
r&�t����3��ө����0���o��
>��ŕA'��T�jO���>�η�]���U��m<�_ZEB���n�Kܴ�"�� �aﴫ&�jJ��މ�v�l���ݙ��x�Y�+�6s!��>7�k���^��}E������+������[-�t4��tQ~G�GuQ5b@���Y�����;UƮ�ɹJ�y�����Ի�Ei�Ѹ��v�#�3��z�ȧ���0$k\CIܒ���1*�W�hדF�g�hrq�N	� /��:��`5�=�CT���!��Q�I��X�O�LSY�����Zhtr�'(���I��9�g�T�:|.�(}.�tJ��N��祖�g*⩟,~��gMn���i*��a��~8j�u��t膁���%�;�ZQ���>���s�>��TY�ʼ�v-6M�M�5��t{;��=�ؽ���>��aH��$GiZ�TV�C���KC^��y�2H��ܯW�"H�3�gQ[�!��/9��TL�|X1��H�=���9}�8\�ޒ�,Rya�����b4n.�	�CŃs�;����>s�-�@�^���2��v��YN�.�{d�|��m
+l7m��{�ᘍ&�j���Ǌ�;)q1<���;wA,*Q�%������bȻ'I/��^���w�L�@� 9�6Q%�͔����Џ�Nw߿3��\���]������}�w��K�!�>Γf:o`N���'D15I���,t���-)`6i��B'���ǳ>���?w�ն+lW򄮫�&�1���Q�	�3�p���;9S�m��M����mր�'SAE�<*:���$%� ���8����m_[��(˟�>û;q�	{�d��%&�����O0�#�Dpۋd%e�YR��S�Qd�}�8ja�qLm�|���L��Q3L2k+�\Ko����R�=�U�c�A�e����lġow~TT�E�㾘Fx]3�_nVd��PHx���V����'U���$�4E���0����]Q�A!�5}\L^�n�@��������a}�ϨN�p�}����	]� +J�\}����m*�����d�L:�:�)/Q�12��|�s�'���g�s�7��E��c�=���Ϛ��W�}�?-9%���:��T#;��h�zz�_�:K���h"���^�}�7\�5Fn{�x_���J�(e:+�-R�I��e>�a�)5\QU�M��v\��>�[*Ԫ�^ d��T�W�^H�(@~��|+���oe����}�ͱ��xa�؞����c��X4H�*6��T�<�� =Kw�^����|jE1�����gO�@!���_jK�kLD!�jw�Yc�MloM�W��m����s��^x��;�P#�μ^����N��aO��r~���w�K_�8
djB��Sk-�<�=,��~�K��&�vfc��5��U�:�
w�61�5��y'������`������QUO�C�al�/�m&t�G���x�J�+|���`I&eo�Ͻc��H<��ʷ:�H?L�j�NVx%I�|	�jJ�ZK������f�̢t���r��4��64P0ˑ�9l^xq�Lo��\c�HNPn<k�����{����Ť�f"��],q_b:�M��)�
|����a��aVW���qe�]��<�-�S����%���������j�g�
?p��S�ފ��B�+e�7J�?���<_JF�u�c�6Ka��=��$��S��~�.n@Wp%��gNN���*3r��|�Zȵ�1��=���nvK��K�AYbd�A18x��K]��Ix��if�B�p,���w3K� �h��<��3�Rd��A~��Kt�3C�B%x(��X���`�^M|}<+ ���J�(�Zlw��)ͩ�M#��}���y_�P0�9?4�=g��"Ӝ�t�����Q�f�N�l�����ė+K`o4��EW�{�����H�� W��Gd	k��?�CO!���1��zt��ϼ�$�D�����ѡ8����n���Y#S%I��+�+��ysI�JҖ���U�3�;r�
���B{�}X��2%����b䝣Y0�,�M�aLP*�C)��-[$q���[揎��9�]X8G�Ն�w��,��e�k+��ڢ&$Pռ6ۧ{�~C6�>,8�^�_Ϟ���b� �W�)���j��~,t��q���B|��S�V��ҫ��FY}\9A)���'��g���^k�v2My)����`�&�����2A��7�9�*k0)">�&��KY�>�v�n3�'v�<$<����dw1{3�\��_�KQ	4�ޘ��M�ޘ+p�oJB��UJ���8��ɕ����t�JW�GC��p����<��]?E�q�c�'@�Rt�"���H�۱i�D(�N����/U��\[��y�B���֜��Ѳ��8jpb����K���>+��J�箻xlg�^�Ӈ�Q��5��R���EJ	��"�j����o�)Ooq���|LDÈ���˛}ZO��U�f�~(�E���*, 3��6[�o�����/�����a���ͫƦ26�H�}W��6���nD�M\�yt$v c%	�G�I��?Tb+Yb��=�۳Og�[�[���=���C��P�f�u)	0(�a{�G��w"t�?�	�;#�ly���X�~T?�FS0ǁ5c�ώ�Ѵ|����G�(��؛):"e�����+�P�0{�Q�ݯ{)6e	i���'�����s�c�@9�1��UIp�ݮ�+z+�)a���7��e�HӺ��N��VS3A���� ���l�9�H<�n�T(`M�kd��[�mc>J���@�nU)ģ1�D���[�����Qz��?�"�UWq�]Y.���� 6-$̌s�y ��&l�t��'�d��d���*���<�r.\ niT���ރ���{�v/E-_ۜ�|zț�³'��sz�|Zȏ�a�59�ͼ�-ȰV�mY~�������e��d���5�+4���vDTK��6��q���@d��H�wK����w�M��݅jC8h�3o9�/�_��Di��=A���r7�?�~��Q�~����\r�<�T��=*�VbQ�﯇L5���@�y��K������ ��&Q蝥�橡�-�4$�Z���T�}Lp�����;P+Ϗ�<�����{�(Q���t���ק/�k�@��=����v�1s���j!����K�_����,�+1C�g��7���?���{V4�U�����R�rS�����ɅO���Q��$��ӚR�&�ƅK��� �,���q�B�ևbA��%Nv��8"�^����#Wb��r�PL�a�JjII�2��~�y�e�̒�ow���d�0�*�2霯v_��v	�A���+A� ŌNb#,f�W�[���0�ѽ8�;G>�9g�G������,^�I��EZ�i�oYhA�rܑtI��>�7�V8���[��a�D���14�>E��Xd
���Ύ0��Y�ud�yR�6lb~]��t�H7T}��;��f��i�_�2��$1i��/YX�U����8����*��Eٙ, P$�D�˻0����{Svw�Hj3��4��P5}��"3�5��,�U����v�@���)�Em�
��ϒ��VtP����D��8�N�����ށ�~Z�*T�;m��!E�]��ȯE�I�g擟��|��ܴ�'/i@[)��F�S��̳���|�u��S�53��s]V{zgIdU�v�(C�=��*���4^�">��	�P�`�M��[?���},a��T�I*��á���-9�Ê'�\5[��c0�Z\6��!�����C�+��M����܋�`0�v�6�wst�p徥4Yr׌��J�6��m*�[N�B�;l�Ì��P�s��W� 6k�:k�5&&J��mگt�+	�E�S!���{�}�Ͼd�>[^7���������`P��#�PKO�[H~}�@�(!�>ܱ*���f�@~e)l����,�L1�ޛ����y�K!� �0t�ɨP!�fǭ<[k"+p�o�;�է�ln�7�(���xDنތ� ��V�8*�j���9p��Y����q]1 ���aY��qn���%�C�N��(8��f>Λ"��1
��=��Xyw}�G�^�WҔ�fe֓U��Jo�b�^ל�'�cy�>޽�cF[^��]ScP�Ǔ�Z�O�I�"E=�̯�~���.�רf#��k���xT�7���BRdq_N����/#���o����W���(�1m�Z��o^�~��� �Op!5�5��6r��=��$\�J݋���^=IshY�P���(�N����/���5�C@�����
�9����s3-�H-|���4�N��.­�ਪ�w�)H�/ ΃�߼�����ٛ��_��q�q�{�Wr !x�.>:���/��x<`;�TQUB�\���'�}��*��C�������!�S!'��v�cve�}��yb�[l��bK8}k`Ʒκ3�n��j�9z��Hҧ=Q�H0��7��Q�������MӣMT%*�����0w�bV^Y�I��7E��m���iz5N
�绿��[l�Nڋ�F��9�IZf��Ws`�AXkD�	9/�IG ���қ����\1n�}����x��n�1�{�O�
P٫�LF���/'g؅/(C'JRl�>M�B�<d;�(�F�����FO,wj� �>����VR�/�?�E��v�4���@�s�������Un� ˂��� ^��b����6361˿���^V���]��z�JA��t��$��7�5�fSTF��f�޸*h�����5��;�Y�1&��=�/^%��h�*���9׆N�
uޥ�H�WNj�R\�J�-����~��8���r�)n��R�Pi���ߦ)�l�6g�qm!�~_fZ��\Y�)|b�����u���%-湐�d�/� i�$�w (�a"��1�����(�VN��W�ϭ)g�Oz��!_ߟ:t�Y����K��^���#�o�P_�P'�������1m�ؑ ���g��y�����_�X���㘋p�i��ދ��ɔ]�[�Ξ���%P,�A���N�]���lL�;���	�Lb�8�	�	h3"],�g�A2��/V�肞�����#Y9%��Wnϋ���6���ʇ��U8��\10��?�)��	�����S9*�� ����Lȁs�.1�kȊA�ӎ:U�����ٶS�V����P�_(0\Y�qa�i��7H�H�F�"A���۵���@���k�3���	���]���Jl������l�9��̏�p���W]��"S�}[i���oQ&�>z�?vZ�7mmk����'�Bvk_]���.@�aa�ِM��r,���E�f���6*���β�`M�sgQ��n�}Ҝ�{�C4�˙^;���dٽ�M�RN�\;>��F�YH�4��*-G"<��EX����̴ܲ#���M)?���Wa���`V���g�O�(�c�@�,'T��mB}���[?��E�\���;�0
IC�>�����������1�I���?A◿��q,xI���F�@7�<�I�(I�n�|�w�۸�J����id�4}�J��Y���t�m��<'��`��:E̎�'���,����d���-:�����ӎVsa\j[�\���x���jg|GYyc�"�ty��|	�{��8� ��58���'��-4=]�BKVDn4Zm��=���sքɄ����<�%�h�ϐ s[MzX�m������:�XP�V,����4�]�@_����E�o$$=�rP~���qm!���+u>[��)����!5ܛ�ŷ��EVu��f'���˙�S��w���E�@�8��w���m�ڍy��|��st$ �]�f�W��'�����sK�-���k�ީ�I�������J�z��"�4xg�� �`��G<q�l��B�<�9Q~��sVQ��?dXr������w��L�'.T*�MRR�ܿo#���
�`�X��N<QD^+��?|}c݁I��K[Ǐ�7|(�L�B���#�}�T�?��R5}\�b�ô w�x��4�],XX�j�C��r^���{�W�e�q	�3��z�i�J���7��dE}v��"O����7@�����w�0���̯���J^Wi��T�b���*T��!��}st��ީ0fy�q+OLҨa���%Bs�N�~�K_�;�V]vE�u�qɛgP���}C���$���F���&���>��ܲ�@��p���c�y+QZB�����o�z ���)���Fa9d�^�Z��IQ�ñ�/���*��������E��T�`ߩ5����aeD���L�N�m}&B]�/=2���6�u�
��W��}�ʦ����T�/��|�.��+O�{���ή��U��sByA]v�k#�������XW3��+����N��܌̮�:���P!��C��5��a�����v�����N^|���&� ����*�wH�F��p���Cjg�����=�;0�CMs%ghuԑ���bcd����HL����L�œ�LB����v{�����=��G�Wu3{����$��c��1����U��_��<	��6�^��a�G���5����W�ߊqw�M9��*T�i��kǩ�y �1�W�7�,�c�t�T��;/�<x ��O4�.o\r&v�H��h�\my�5��~�[�W�L�Oܻ�)����� �|8�9�|��jvI���؛)m7S7ӥ�Z�'�IF�x������e�z�C��>�}��`�}9I%���ì�����o�g�cX3�������ؼé����Ώ�F�[��i���2�+�0$�S�fR�z���B���C�#N���zPa}�l�>��ݽyAXW���QA�_�ek����b�ˆI���+E�T�s^�/��΂�[+��������l�T�kgD�Q�N�]���=a�g��8������fP+�6w6Yo�=�#:mт��<Y��C�'��d�#OR׵�Y�{���6�oe�4I���4|t,��O���*������](�]@��EѬDPCC��J���w�ZK�F�=N8%h�x�;�����o�&l��t���(d휢{��_�*3�~�֪HUPFC[�`���g��b�7�g�<P��u�ɡv����գ�Ϭ>'$�-�x��[`��f�U�����u�ހ���Hl�!t�!k��,8`ݎ����}���W1�N(�oM�&	�|���j��\�2��iw�2�F��B��@1�۝'I���v�;N<	}-�t;.N\�^��{cA���D	��\�8�\�?�K�]Eΐ��A����e���W7)k�s`cY�ޤTR��{;�($����v�Kb�:@.jd�Pwy���$�k9e���f6s8Sa��|���t�=O ���G ���_�$�gKO
1�.^ů��Xe8iHn�|��8��]o�Ն���)��@|����ξ�><gt�L?�S@^ʔY�aT`A니n<�P��*��>�E`̱�̵�	m�2t85	��x�^Zcz ��f)
L�1���*��m���Z��9�i��!n���H4�y.��� ����'�6YD��p�G�\�X�RNI/𵪯%�Nۿ`�-���� ����:V~U���x3w�m!r[��F���eRoL�����(t�JK�m�9�M�2�@�]������	b��5I���{a�y����!��c���j��cD�@�x�����k�;�{K:2��,�"_���D�J��y��AI
E��vቮŨ"uN�`�u>�oi�F�C�~���Ӕi�&�@C��ʏ��s�T�j#��s�dK�j�n+��e��#���zo�?�=��ⅴ=x��	Gᩳ_�f(|-���|?��׮�OJ�ԛ���Wљ�$ql(�I�x��&\u�#�|�i�'jsP�y����rydXO�`���'�_���'�_�3r7�x�䶢W�K����l�5�ȁo����6:&2.���K�������V�ho���Sc=�_��Iݐ�J��Gq�������˳#!N�#,����|�O�ؠ�88�h�z?'L��`���):K��G�n�c����n��";�U�
6��=�c�o0Xlf<//%��;�}���l�ʙ鿘��å��-;��̔�2;gl��776ZD�3@7��y�Z%���)�ӓ�3��		���5_��@U}�~�r۱f��V䱪o�pedzq�2k�t85�=ԓ���T�l'��6ϳo n}������,�s�,H��_�n�̊.�8���q��7�-����Ƙ�l�wta�5ke-�P��\3�U�$�" h#P�n'��`��x��aM��{55gX{�C���N�v�UM�.�Jt&������-���#�E�x�\��\��5�B�֞�s���7���H�Ū�X$4J��B��dU8#:Mi�а�7��5Oua�^�5%���o$��3�$�$�v��� ��$m2�Ag0[a=-܄�ڝӰ�~\�+ `~��^���_4п�+�<Elq��s�@�^�3^j�k�����`'F)0�à bNAŽ���!Ry�A���=�q%xsʁN.����J����n��~�����G&&�� �F�x,	^j��5���8��Vީ�>�I���`��\��-� e��'�҂?�u��20�t���\���t%q���Q�2�,0�+��!��=P��Xn��:��Uo�����m�3��u5����3�֔�ʩ+!�������+�ak{5����sѻ6�St��mo,b�Cy_@n��vc�3tc�b���z[����t������Gb4�P����k�W�����[���Rn:���$�S�kH�*�víb7� ��g�L��𢕺�w���g?�����7��(���6�U]���Q.m��1t��
Ы\0���4�?%;Rd*21w�ܘ�u��|tC�= �pb��Q���C� �c���ێ��f(\Z�~��O*�Mn���l�3v^�C��������L�+y�21��>�:�Ƭ�<ۗ/��pW��2�� .��G�}7�l��#���/@)F<����4��}�(q���Ϻ��"h�7�57j:o"���ᖭݐ[���5��u��c���c�t���,)�����K:��̕��K�L���G?�j�v
����"�V��P�6��Nc�Q��Ӓ�)�W��vp��L���W#���#b�I����Ine"�Xx��n�?M5=��p~�����ۏf���S&l�qqz%����t�=�?��ϑ=��ӟ�U۷�E�c�� +�d�������?,'�U�I(��	w:̞����x��IUZ7�I���j�"l�|��:��7�}�����U�i���d#����
u���08����xh�$,/����(�7H�m��08���m�)��Z�2�J�Q��>�.yL��R��`�7���m�~إ�W�v���ji�I�-����ED5Mg���Z�=?���^lټ���^�n�%��$[
�����t�t>w�ܽ�92�E�П�;�'uʃ{5t5��&��h>U��6ew�go�\�]��SA\8N�=�mL��S�`up�[qO�W��R��Sd��N�h<Rd�o�w�k"�b�y�8ʫ�\�VH�C��*��Y��a����/���v��u���L�#N�W�L|  Q쀱�����g�:E�^�w�|��&/W^("�Â�|��W;��b�ѳ�A��'��<2���q���}��C�`�ۥ���SOEx��M�"ɼ��_�i�� 0sm�ă`��sx�a�I���G6�^��=�to���}��wz��GG+^�!�����J����".A�Q���R�m�n�8�-�y�.\�  ��C�U�b�k�"��]��V���m-r]�H��B��[b�̐65�ae�%���]��=|���#+���%�.��,$���3�Z?��e�i���Q��xR�ȃK#�� �GMg���f8ki}RI�ɂ�Rӎ�˸�������Gk�c�8�OH1%:���A�{�W��rt�а44,�+�2@C)^;ӓ����l>��^�j�b§�
�:�O֓=m9�5y ��U����Q��
���#�`�f�����V+f�f�r��2.X�ΪCu�<��x�7�"b��������B'C�҂弯9�?��o�Ȳ�6Pv�	�p$j��2�˓���Um[�l߼+T7.d�N�^Y��~ 2�.��Sx?��hm�7���˞�6��e���["����F@�v'LA)�Q�xp����0~�T��5�ɯ1 �m�� �V},�~�o2��1�t���E��rI*��ێ�КgY�}y���Sr �.��@w����P�� )K �,�iCj�sG�򡸭"�(؜+�.�;չf��b�S�?��I�zJ��7��3M�Eak���Y"����wϓXQo|9hRM��[��gW���d�R A�](�}z`�V�F�r����ƫ%����{4��l�Ǹ����m����b���ۤ@�;���_)*�'�N0G�m>繥���C&lώ\E~�i�6B�#fXb�g�p�w;2�5�-�.�l��T ]^��狌����O��!�M@{�[A�qw��u�{nZd5al�L{v%��Č���
_�6��D���f��K�g�uGmx��˲��CW,��R�!����:��`�p?Q�����@���B�,3��w��U��*�n�^��cM�.G � HT�Ұ�5i����3���/�gPu�3�թ�Bf{&_���r�u|AÃ���SJ&��ĵ���|Q�:��k��X�4��Z�~݌����)�h���~����gP#��@��/y������)c�"��s
���p�4=�����ƞ���~W�����T�� q�%��5�m�ϭ�,T� ��=E��g��cq�=G�
Ё��Mk-.�,�&��ѭm�Tl�Ӫ��ye�6J.�� �?Nu�WzXf�N���=��������o�_J�l�W�;Y���ii�-��]���c ��/��GmJ��j��"�!�5X����T�`bF�d��A�R �p�m�b��牋����w:D������곘�_�k�����;� �����7��.����M� RF��g����i�V=�rV
�VbY5��K�:8)B���/��Mw0��o��kiAx^��B�@{������/����T<z~���s��H/��1{'������vs_N> +�=~�v��f>m�w���>�֏���g�{����M�����Z����M!������y��gK����q�Z53��q��Ǝ�����:Ig�e^)��8ڱ����=T���f� b����;�L2�������ћ(�87�{6���&������&��<N��'< �1�����`�[[U�ɸ���YC����is�ZC+�B��~����d���x�����r��A�ϙ;��ȧ�A�me����y�oƳ��2B���RT���>%O:_l�6�;k1;M�Aڈ�t�9�赉��Y�3�VV�=u�&kT��W���5&ژ�^����M��TZ-'�Z����?k 541ԍ��U��*d)Y�)�zj�/V\c!	��s>� x�40�Va'���v+���C¯����c-&@�#Վ_<	1���&I%|����z>�z��hG-<�ѿܙ+�VD�bف/T�U�;�|E���&�xoޥ9��Zh��q�UM��Z����.qm�u8���=*����NY�L451Sc�k|�tLam��EeŢ�w(@B�S�z���ݘ���<�н�6�e���=�E��.r��)7cE�*��5��u��ށ��*+�l�{ߦ$������$Q�akE�J+կ�������+�+$O��N������˹�^
�����#pk�������?�s�;���G�I`�6� ��'2�!�׺�[n������taH>�����ه I�% ��!��5/榕��l�t0<�����Y�@�!��8�Q���Y�>l\#�2r�;#��_�\�y��F�|��?�T(�|�Jc(|"ek(�������
�&."���,dq��_�Z��������e���Σ�����d�,�&ɀ�^�F/�Aփ����j�w��$[��5���h�k�Q�5��#����>R��Y���"����D�ʼ�{�z�`��䧸��S�WB���;>3s�k����_qmT��uF��� ������4�7J�S������������{����u���W�v�q�XC0��m�1��ǵX~�3|�����폥/�ʹ���1��!CV�5�B����·UA���t���ND⃶��fR{��/�ie�/���ʰ�q"/����hKn�����v}�Ư��U|�Л3]� ط*w�5Kf{?;��@0H\Kr~�A��N��"9+�-������ߢ8������޿���O��At|pDD��f���'���.��.@r��O:��_�堳2)g�9�,�v|#�zl�2h.`�5���S����D���od�8����K~h�۟5�}j��J_ �������5�Nf��\�����_Cg��e�����N�2i?�_�_�]��Lm��Im�I0�;�f�-z����ZW[ID�(dd�'�r��� $g�߅tˇ��[���uЉB9;�^k7�
��Vi��\{�����{都�.|43~��Q��"HwA��F�*(H�ދ�( m��! -�^�ނ�@�QZ��=%����?�_w�u��Yk<9���.�~�~ߜsR0{��>]�O���*���9'W�E�U���6#�#�E �Z��y�tj��IEN�G�~�s[��?�f��Ku���{�t��o�A�"��,��D�B'y��rƉ�ݾ�ވ�j�g�U���r����#�A�����_�R�i�Fq�s����Ŭ�(�\���!r�O��ǚRW�98Lk��� ��KL�AP֔�y�}��a��\�~yQ�3t��-)�Ϟ���_42o�'��-B8u���8g�@Z��D�N~�*���qЃ�Frt�A9��R�n+�#d�����oE쓧Y8ߪ����8Fg�,��<��Skd��p�WS��r�����k�f~�	�����{+��&'�����h3��.���Hea�p_$�B!♂���rY�vS},�QD��!��i,T��:H=�nչF��U��6WG�~��H�ͱ��Vϼ"�9��YcN?���:���x �l%Dy[g��F����r�g?0#�>�ꭔ�'��1f�ӛ���j+��=̡��da˫���{�Ǉw�'!��D��5�)��Q`dY}�?��Qn���C�"���  �1��8 y��i����۸`c:�s���a���K2�:(5]����יQ�5|V�oKa|��K	u@\YZ�M���G�)�����|H�m�T_OW�mݿ�+5�Jҋ�sx�r�!�ʟ�R��u����v׼b4�5��tF��c�5F��)H�8ʪ�V�̖�U6n(���Ӹ�-ڧ~�? kU�i���b�"�2�_v��n���?��'��ʟ+���2Dq��o;�G{��)ɮ���Z���G��&Wȭ�#Pfl��*j��xO�b���G,�
Jl�)��Y6����;Q�W)�^=ao�I|i	�D���ҩX,��E!9n��g1��l�]`d�zPV��Ā��*��F���k��`A� .��%���zf>I��)V�5�ȟd7�n 
%k-��BI�#�B��fx"1Ů$J����@�c���B�mwM�	x,�qq�m��u0;��˥�N��9�2͐��YͳTV|��T��,z�\d*v y��wg�{E����׈U�D�OW����
4�/�o���@V��$�{�*FmY�r�Uv���pZJ;���#����}�jH+��U�����:.(�I�䷪o1'�3hUt$F�۷�I�3Tؖ5B�K���/b�]�g�/�B��~�|WF��)��;�`e��y�%���0iw�IĊ��� �͙���ѣ�X]�uM�IS~&�Gtw�g�N�	�Ո<vK>IL�pn��>8�z�։���"�o�UYU��S	��o��)�L�Y�W���t/}�>�=C�@`}@�� ��dv��t��s��_1+W�Re3J�>_F��8��4Q
���o	�F�O-��FFc�zF1�ԗ��x�u�݉	�SԽg��	�jE�S,�?��t	=�򕉚��fz�ߌ+7��߻ᗃ,�,hyfT��Y���,p�r*��3�]g: ���G&NIBn1�VÞp�������4��$~���rU���G-�29�{�\3�8�J5�k�a{)̊�r�^.j�.x����J���8F�tX�"���� ��$u����$�� ���I��x�+W�Ӕ���.���� z>��ܾ���<���#�
\+7'>����Ox�w�]�߼����~�B�����f����8)�S��r#3�V<{�۱R��t�KÊ�����YNn�g={��9�KUB�c���{�G�G�Y�H���ouM�� Y(�^Vڃ+�q���oZo�c��=�Q�.�jԛd)���H#$��	r�#�l�$�"{\��5*2dX�����U������|��?{�f��
`'�lN�9�r$�0�m��҅�$;�r��=��0ҺY�aeuLo��&Y1!n��)�s�W��tS��>!��	.&>~v�1��+�?P�K�Q��{�얺�u��SV3ho틍y�#-a��>��*�V���@vm��L/M+��@�Sr�Kesk307;F�W�>��������Bkc�}�����E]ԒӸ�Cg,3����v��1�q�����3+~�*�Q�{Z�]�~Yh�����w�!��&���֬�(@ղ�'VzJ�e�K@H��@_���Oֺ�Oo�e�I��avT�����(����_��WE�,�)���ԟ�v���?y]]���v�[=���7�Z����o��U�,�+Z����;~��~pk�peeWNˤ�tk�.�����8�+q�3po�����.{�J�a�v� �� �#���tWxzv�54�B98���m�"U�W\C�@��^��1/CW�i5c����S1�}����Y�	�J ���.ӿ*2��:�����s�q�х<��)�l73�,pK�p�+���c��R]�{���3���w��K[��T���k��KՊP�LMWsC=;���s}���i�tl� �&7����q�c�g����Q�l�y�g_�K�^-�������`������m��wW�k�r��e/�U7ơ|���O��S�o/w6٦���|�Q�n�飧�*��T��aq>S�,�";J�k���-�ǎp�_c ����ےd������F��"w�s��<!�!���8���W_��Ԍ�xδ6V��E��=o27s;��V��B�A����G���U��*:HSz10�H3@�nlՆa�	h]ɍ!�mک��&kooKY�|8VF`;�*��H�������%��`p�'Ǘoh��^Ff�&����`�{���[;%X�Gܒ�.:_2�^��2��u�9H`��'	�<�C]ɽw-Q��i�� �k�����+g[�B�S���Wf��	��+�8H܍I��.⣳�ՉE.6�O��;/ϕ����Z<|�{���ڢD[�/�y�>�c:ut���RǊ�����j=	g���0��X[$/�O�j ����������
�����b�$7b��4�2��ţ�X��b�v�d�z��'�j�H���T+�@�o�7��"r��H���ys��$6g���eO5S�/�a�X2ʗ�I��dU��b�,��x�b�hF�Y֞�"�K/K|	�5�K	*vb�K؈�����^����o��lx˄�_-N �}�q�	���0I3�9�S|w�n��<��뜅邻 ��e%M���jG�ṡ�[O} ��Xg������m
���(ɝ;,?`�-B򐔧�xT�� U^$oa(N@B�_���b��zCA��^%b��-������w��J��K�-� �TV
�6jƃ��)�Ȱ��fc+�Aޱ��q\��_�.�kg*$2���ܖ:q롷�(?���󀊖��E�d^��=���(��F�׺������.X���l�Z�=�t��"�5L���{�oS��+�o@��v8��X�2��DUZ��K��x����K+��j����b<)~���<-�'^f���s˝���G8H�ɟ�����֤`���`�Z���|�;�^�hF�۩k��[N�	�\Tϧ�|���yϏ��gGqdl�\���bm!�Vda� ���O�j�8@�֫����=�*�u�R̍@��y`�&�����p�*���k��`w���p�jk�>�"Sġf�@7>*[̿��a^Ü��޽Ԟ���^�o`P�t�ʊ����W�+<���1_��}�7Fy�J#� ���Ү֝�O�;�I���,�[[�؝&��ƛ���̷;�Ag��D��admQ7����&%���x�8��qL�v7Bq�n�#�H���c{�uA��0�� $"��v	�fI�[�T9�6^�:�~����~F �3��Kx�ȈDh@�)"���<���SMd}%N�kn>X����g 5}�+W����Rܜ�����v}}�����֕Sl9 	&K��O���C$�+��k�_�dv��ZP�V��}�n��Ħr���P���:�sR'�g��i= �"���J��{9�0��_�,����^qu���-��B�y��W�UX��S��� 
��6�}�~Q�TЍ�5sn0Y��07D�O�e��P��'�v�&�H��.��f���7�3x���<m�n�`�1_KE�Y@�����$�T3�mGB7����/{��u}�pMD��)����+�Z����x����!�(�:��@���Op�¿� T%ɼ��[_M��� �
LT�l]#.��6��6bv�R=�?X�|�0r��+�� b��������zS�(�k�%5H�ۡ�i�����2�C�KK�+l`�IRTT�0gt�����ػ~���ot4A���pQ��?�@h�Pcִ��[����t�b��������3cAlxF��i�l��#��B/fB��J����;H�-..FAij�ɐ�@��е�$G���-z��tj�E`n�]^x�b@�)\PPi�Ę$��x㨈z]�
!A��{�[mv|n/�3�rm&��u�����C�N䕑�g6�U��n��Cg�6ϕK���j��ޢm���o�3�-Sɡ���9Bl+�K9���2��¨�h^���*�5��V������n��0i3]
��=M'�����'!͟�)ߒ�J�j	�
o�:6���>R�� !Įnq>`{9H!Դj|o]M_�>�m-��N#YJpr~ZoD���zO1�s�g��_+=���^���qvވ�&���)�}�ͫQtp������n(V:�r#�k�_;��g�������T��S	�v�����C�4pa^/YUU����!�SnÕ���m�h��+={��+��H�C�L�3q��p7R�btX��pKt�y ��D#P�_�9��e����ˠ[��w��+�/҇5�&t��Y�농g�O�UK�Totуޘx�v�1��m��|���*{;�����RN�u5��S�LU±o���9E�Y���V��٘2,j�����1��!�1y|V!��I����z�|U[�G��7�͜;�g� Ă(���m~��t���ݾ�<ohlh4�w�ٕ	�5F�'�>�䊬�oo�3��U��ʣf��:��|"�rdׯ�	]cN�nq����3�UܲE܁q$s��׼�� �G��t���$�;�lT�1֯rZ��3�"T��S���z˙�n�7���~��)P��F*�������z!��#��C��G�z"Q�a���R]�m��:��-+#I��Kń�g�Y|9��Α>M/�\�\XR��� ��s��R�&���w􆉣��3��Q�2��@O#��-���I�-�ܫ�4�֔fsȧ�'��ax)�0`*D��x����^b��7B,�g��l��D/t��Vk~d���E�3����7X�-NUpj�o4��G�2
' OK��{��1��5�������P�}���\o�zn�z#��/JA~��a��kIto�+虚K}��Qg��݆���9��u��7�֗A��;7��7h��s�܊4azl+�Ѻ�/���f"�f�y4��hPE�@+:\Z���7k�!0X���F��$��b._U_���Y�p�JHk�����0�%ZH��Y���r1Q>�3���@�:��3Hf�.�NvHc��/O�D�8EÁv���ߗ!A�������#c����0�!�S�H�@�
�2�䢇���bE��0&s�x���_�l۽�3}���﹑7�#�c}��s������wC"�J������z��[-���A�g�`p�`��2L�>��������,�p!H�/��"�;+��-�$6`4���wD��jj��1�+�J�m]��iy^�QJ��}�c�9:�,��kjC,�2��Gn����V%���i�Í8�N�׍�;�V�B̜��T��=}:��RbފdT}������Ky2���P~� �F}b�zI⢝��b����"xiW��FmU A�����\�W�J_���-De�ˬ�+�u_���q�T8G'��M����J�։ !�K�!���FE�+���my����1�Ӆ*w!��i���,H�	�>���z���u�^�zc�Y�ż���g���n�us��ZGsWY�	m�Qm�n�hTp�a��o���wCu�Qs=y����@k!(XE9��~�ss�PHz\&/�{���m���C]T�{V	�\R-sƱ=P�'��w`5���|���y�_���B��M˛p�0��l�a��V����8�=�����M��n�De�@�Ǐ`󆧌��Oon�{�s Ȕ�r����/r��P�WCȌ����4������Ό�������QG�_��NȘ�8a�'{�v/��%P���F۞��+�0��i�}U�0��z��x�����mC�� �ăN�q8K����v����1˽���D����|��̈́K�P���w�'�% S�w��CVJݯ������7���/�+y&�����k�y�X_Uܢ?@s_� t��]�_f\u�Զ�Si��L/����q'�5>���D鍻y����@/˥1��'Ry�|9��r�α���264v�48J�ɽ�g���o�*���vns;�2�:��e���- ���x�wo�a�Ҍ�ǃ_�H��j���Xy]��o]�W�>w���z��}�07竐�6�6��]��.b8�nl��|�m�:$��6-����^�o�N��ꘌ��_!�8BL�w~��k�el���N�v����I�yE3��7��n#7�{t-�z|�ɯ��Ef����CU~�7ꣃ��� w�H��"�^l=ȇIf��Աl]#*?�t�p�5��lҘ�#�8�ߴ�9�Խ����=��� ��'�1/#�{�q=������j�K��+vt�;��À���}׼�ja�Ѐ$s؆�|��=��Ώ�_��6��sx&��Eu�ӯ�/8j^��]/�ڸUW���s�j�vz}r�6L_���q7$�-<Ȝ��s��xQ�yH3�Xܘ�ĵ*Q�y;���6����6�/�B8�1z�"Wc�YQ�k�4q����H��w@<��f������1�1�����c9�}�
��Y&�F�@�y�ck",+!G��.�&C�÷lw���K<��x�l������;�贈�V� ���-\���k�~:䎝䁈%G�P���,�N�k����ޞ�.�0���%�undf��dn]��a�Y�g`���܋���>� mb��8cl�A��~������;�o�/�&�jx�6�]�] Uj:�~�]6IL�"��9魕��M�J�Qq�.�n�*R��e�|�3u�Vi�s����K�Y!�m�D ��[u��$��7����'�.o���F��*�ް����Sޡ����	���1�����N� �W�=/8���إ$���%�
�G��4Qf�A�Q�՛B���E7�r[<���fm�.?��������{�|���IN{IgU�f��%_�d�s�jG�w�0��������S�+OA�O9q��q��G�Sϴ1�4On��7���M�j�� ��x�TJ�[���&�<G��~���
d4�3cX��� �Ȇ�z<�LUL�&b�������W�hX䖔!6��{�{T�~mÆ��>j�0����r�_�"�(���I�fO�2 �z_!@NW�}��q�_>������~��O3����y�ȷ>i���6��e�9�V��)����
n�*�h ��̍��&G��>Fa!S��/~4@��n��9G[>��/�xz���ӹa����?�1�Z�B���BzC̤,��������S@R��&ō>��]N�
��g��ٚ�j��F�tGo��*�f���j�xׄ#0+��ж�m��zȤ�V�2R��k��=X���?��X� �E�/^�{^�iqQVD�d{�?��n�����cS�U`[����RĤ�S ��TR��8�����'$(��X�"Xok���u}�D�����\�,bp��h�A����@hй�����0������]����h����Y�X�_����Ӣ@�X�rX$�x���%��c�XԓUOeL,G��-cօ��Z���(�	3Z����~�����v����V�3���@���0$(�X��_\�Z���}T��﷫��G: �a^��$���F~B�g��m`Dٌ�N[w�<?_������m"�\�q	׀>�g��z��O��3�'���
��s+�Iw����QT��P@c�� �_�}���@�h�g����|"}}|��i��0t���" ,DH�vC�ר���k���:��Æ=7ȮPle&�L�*ف
u�����RX݀��z�����β��>;�@�)�:�l��XK�������N�:gC��`1�5����
u�;c�#� �1}9�U���~h׫�6���Z��������f<����c�[g�i�0$�-,��ĵ�Ny���zR'�4�Fݎ��� Z
��\�G�$!Ɛ������-�p�� ��J1&Zz�/Vzz���ֿ�X���]T�-���/����l��sk,��D^����x�ǟ�3�K�^��N�;�x-���os�sq������g��-d���W�y�1�rY��e��	L����fW�&���!{��w7[�\QU6��]�@�^�s����ƞd#��R> 㤷Q�e�����
!�(����	�)}2g���!Q#��C�c����X\E���Q�h�������5��kR1cvc�e�� ��C͹Ț*��N�-AX�I)�cs��*�ƈ��P�Y⑪�Y�#��+��tga�j�[z�2������;oA�DM�Jc��4y���V��cJ�O�C��[ ^]���U�;���8�6GX��;�&����$�H�Ϳ�y#��b����t�e�b"�탠�P��bn�ǌ�x��X�7��yW�)��=��=�˭ixP�-�T��L�閧i�G�d���6I�67�� �o�nxb�t�����I�6FY���l,�=4';n,�`��w��_�U�+%�Bum�m�o����=�#�b��노�"j��\�)�'t����k��O�&=�f���@tq�YB_���w�K?8{�v*cF���gq�!j��eg��<���D�\�����3	|ԏ,}���r������p������k'K'Y�5�\G4�KՃFF�d�"!J�j5n_���V�]FS�����l�����>����hw�Ul����k_�Ұ!����w����)v�G�v�� ��HN����2��:�8NK\1�gU&ħ���I��L珙�#|�~`#��򄇮�θ���9$PTB���H���eU��E�jם���[ë���1W�_��^}�m�D�._H&���)�I]���݊M�`��K�J�+#d�W�^������@�ę�lժ-�u�~�iy�nk�w���W�'V�OGlW���[�5`���d牶jhO������XD�� ����;��rQÿw����MN�\����*�K�A ؽ������yF�yɮ�0�	11-��?����!�W_�����m�f�cϘ�y�r��?d��[���7O 
�C��`�_i��Ǝ:fo�*ҝմĺ^��cc�=b��J�����!��e)�t�c8w*Q��d2�HT #2i��9�zȫ̲Z�'#%C��*���ٮ��8[X�*�T�_�p!�2��^�I������ٟ���>h�����������ܵ�MJ�~���Y�㐴��Rl���H�4A*��t}a�����9�Uy��]��e��o��%�U/����vi���5����i����Y2�'��C-�S	T����\�)�A��tS}��ݱ�;�`uu���li�Ets�]��x@�j^9o�.o�D��ƪ>��,�|��,ż��'�m��&g�#g���XL���R���S��� �:��)�a���o�@�����j���6�4�R���w�;�AJ�4�@��&��6�98��E	��4��f��H�ʉ�PI��R$���W\5�ζ�	�؍U��z}D�K��ꡆX�-6s4g�b�mb���.Q�6ѷd:̵��dT��O��xɼ�,6l�-��͏�p �vM�F��a�cņ�0�����s�`�E6�ա�\�X�/�zyM��j��Ʈ�TE��ϙ��|y��+�ٮ�����1�N��F�}2�n&B�"��t��D���l1ks�Ғ�T��5
6���C$�1*0b�3���np����̋X͋{"�(��<��P�� ��e�����Uk����I�,�t35^�_��U(Y����/]ƃ�FË�y����fG�=*��8��Ƴ0���5T4�y���� l�*���X�X�]Qܽ�:,,e՟Ӓ��M7[w�	!�a(���/o����\�Y�u�x��J�i<T{aۗD`��3�DW������r�=ҕR��[\��CSyR�ƺ¬�t��+�}�Xgn��䎱�Θ����0��hv�Hh��[��ޅ�����Ǭ�;�n��Z�����R�-�М�)o{��'�)���kLJ��%]!Zx-߼�Rl�#b�#�:��}���~��Cp܆ +�д��e���fѣF�P�Pj2�^�c1a7;f�&�ی��.�F�i�yvʰS����G:s��Ꭲ�����t~���6V�M���B�Fkqp���C�����B^���E
���zwF�z�}d1�L�.�(�y��x����~�5m�?oT.95��!�D[n�"]#��.7�@"_��}�f�3n��q����X��C\�S��!�@S^G�p��@�#(��z��[�5zn�;�]ݓ��g3���Xm�9����06�~�2e�dAiX��1�w��r�Ň߳����d��<�����7ǨwW��kC�H��U�4/��ʒ^U�8�zw�:��࢛G��vI�j|߷R�x�Q��{��#̽�!.W;D��RgR*���z�e?�b8o4���5��</\�����m��k��a>9�lpw!�z�SP�Fa�n���j�a[��� 1���Qo l�˩�4V7��	P,��V�L��0Ow�f����xԏ�_��oPN��(C��bO�/�	4g6|��Qu�u�¡{l���d���CA�MFv�?�[R�<]h��H��_�\���n�8���:/%P��X[gZ�34=S�c�Q�Va�fr2w�}R�%qaOD�ce��a�n�?��`u=-˷5Rc�x�dو�L����w�	��K�����,w*=�.6��ۮ�Uo�&xb��Ʈ[QU�iO�O߬ߏ��s(f�j�mh/86(˼m9�.o����t�=��C8e��ZԱ¶�B�ٻ���eݹk�:r�wP���쀐}U]�q=��2�� �ePUB�=�,T;#���'Kץ��*ܟ����;쟕�X�>|�-���f�k�|�Y<��|*�|;�u��E�����_'��Y+g�ެ������,>�a�ݺ�{���;�y9rAw��Qd^o���n��ey>Z����h 3v���^$���{�?��W�Vǖmk�9�ʪ������L+��E��d�	�^k+��OV���d�>�~�ˣ���v���y�p(zV�6`�m������O����{�b���BZ�����T�eX�m�+9��]0��J�+�t����Pf��XY6G(u��09�+d+9Y�b�ꄍ�Yloj��a�3���:��������=��d��r�����	���%�:p#/�G��7k��U���S��ݑUO)voB���FJ��it����w�{��{�a�C���~���1����\1��p챫!��g��Q�(9��ȅ���ʬ���v��d������1k���c"�s�±���e�N���կݰq5W�-  ��QNU��jrvB��X���-���������U\�N����bY�e���}���5,��tGxu�Y��Tx�R���S� C�� -h�})����'���~��q���'��q����'ݐF޴{�?�܏�?N�8��䏓���\��B߰���ۍ�^������?�~�8�q����я�G?�~�8�q����я�G?�~����'���Kb��wuU0�����tR�׶+�O�Ҝ�t����'-/�oӇ�'䜫°Hޯ߼�uH�Th��~��%��OWj޲�_�RkP8]� t���W�YUħ+��v����z,��w����[ۨ5�_�~���߻|�����
����5��9���C�?�gK��c+���D;Hl�3����cW�;�[c�E�.<���w��+���.�#Q��P~\ $J����W�=T����D���X��Lm�����?%�1@׼`�9al��Ο[�o
.WP���i.��o�W��R�7ܟ?���25=@�q�',:}2be�V�7�}�p[�T���'Ta�B5w�C�z�tA�o��������ރ�,�'h���E�^�
�>���w����4��ݮ�A��2޷!.**J�������P�F������!�ŕ��r-�2&E�@�qG�{N�w_3�u�J� Xrξd�u3�������t?vѶ�nl�ݿY�٤ؿ����X 3���b)���1]t\��)UƓ}�
�A��p�j���OA�u��ut�����ӄE~7�2v�����oǝ��2l�j�����
�϶���X���4� i�?�]H.yc����Rkʻ���VAl2A�%f����GI'c�<�Pj��nh��G�[E4�"EUuuu��ak�������W���}?{�:;ĕW�P�<�!�"4"Gb߉��)&���s��%<�mM�87���($婉��r'$���L�Mvy�:�w����S!uMfߓ]�����*�M9��=�]
�ː���+㱌��ꎷ�^4��d��J�f�
��+L�tH-��t�20�^���8'At�hk;����q������	�a 	�<j׃���y�o_�%(~&Vk�U�kY����@@�\*	Z::�gXA�֐��z�x��S�����!�V�[O-�Pe�>�9��f�xxx�
������K	��� ���b�)F5_%�o��뉚���:}����5�wzy�i�@�;�������˷wv]W�o]�i7��W�p�:J"�o�Rr�� 3�333P�e�QLy�i�#�5&���8[���v�$t���:�P6��e�/�W��i�+VGԨ4KT�cg!��r�n�	�M�B�{�vή�����H�ґ���X@��(d�����k�uThzH2���L�����]G;nb����:�/�TT� ������\c�cs�(U3���Z5>�+PJ��W� ����a����E�n��r�Q3�e�O)D�\g~~~�<����4�ɡ+$ O��;@Ss�
\��@���~�vUA�]5���7� ��\.��B7��@��<��/{U�Q�~Z"�H3������_ ����s��tv�`��]|���!��?�/W <>svH�fr��xG���:} �j���DӜ�۾��]�j��ffJs�W�ڿ�[5~G�淀�-���PSSs}9�aߡh���ȉY ���D���PSB�\����0����g���a0�q�D��)��./(Xۄ��˚�S#@��8���Y�ͥo� ��i��%�#SG�����02�h<�0 #����q����Xg�DONø���x���%����]�=��!p �>�̖�p�c]7\*.��ߟ���9k4��9�'�XMHF��CT�@N2���@Q\���i�@��@<��~��;6P���Ls�R���%ԣ��ɭ�pӵ�W�A�6 p���B��09�M���Oi�>hb��-U%�EyI��>�f��!��ζT�3��9�c
j}�Ga�V��!�f6�x$=Х��㱫�{w��	�TKO���C&��QB�U��~Ԧ�&%-�����Cb�u۴���IN����$���É!O������V	93KK,�L���O�Q{��W4�
S�{Z�L �� x�WdA��y�WZ`oz�9���A�?x 'X[[[�|O@/<4��z�+M����g�����Th*fȲ18��P�v��A҄��my����n��z������	Oy`��e�N��in�x�wK#jiU"|ͥ����˘�L���Rz,�2�<Oʞ@r��/ W�`[�[�E~0��!/�H�F�("�9)������p�Ҡ�#�b�Ă�oY{�Z�0�}W--�����F�8|��3���c�T5A�Z�]�J،7U��}���0|���$��K�
_n��I�ﶴ�S���+�"�!11`�zW]U���_v�Z�u<�<X`.&x����cN[�s}��<
�4ʶ@�@��`N[`���չ���av���"hN䔑�@�_�ψb��`we���}�U �&|�Y�Fu�W���F�E|�=��^��ȗ�y�@8����pD>�][d�p� v��c��n�#Ǥly��`�lQ{[���
��#���7L��,-�"T�Q�g����Z� ՗�ke���&1��[@mX�<���%�6�$`8�ځ?���#�����d��@�Z��#�}_6Ix
c�%����,""��{�z����j>��- _<&:�8���Q��aa�!�@>���[QV�1�i�3m�EcژP�,3�3�x#cc��Z�u-K���$7P����'����u��m8����aB���f�2b�X���c���c��J�K��[�a#vz�0��ɖ��	���67�Z�sI X�U�A��7B+ġ0�*�2�݉�86m�Y0���Cb��|�Ɋ�.Yba��i���wIu�h#	���4ʹ�`�4�ʰ�P�/����0=�#1� @��n�E�>�e)�D8�\��)�Y�xR��Bf[FO��8S_�&����r�(EV����-�� ����#u�ڄ�S5O�f=Z׈F5�����K��7���H����ճqp�c!T�j�^N�uX)9y芐F�dM-�r.l�Na��5��iJ�4_���0&(�m:�u
5�2�����IE3��f�2�bꞽi4��zD�꾆��iH�	=��c}�
�I�^�4�ޛ.w�!�|���BzG�8���g��D�6+ ڹH��^�Jo����1�)/h�؜<q[���P4dL������n5N4�����
Cm�slQH�H {����v�kceilE/A� �������j�F0��G;��(3��j�a�8�ٙ���r�X��kC/Vk*\�AՈ�	=��G����4O"a�rv�&T?qvޚ�Sߎ�:�1,ú:����>�pqw߽� Ʈ��f]�yI�)%$FĆ���a�L533s���̯��$���@�E|c+
F0�6&�$Z]aUCID��Mڧ݇}�P�|���X��������U�Z.h���A�a���p�s)���C� ���Eh���u�$!"��QR���"
��аk�/� �!�/�v��j^"�F���JX�q��i�z]�*$_zHz&	�	��&&�H����*r#3+�R
���;>��7�c��q�C<u���˦�W�"+���t'��tͯ�3�Q+��Ht� �����+�2��,%�*�J��Vbh�:���=�bʶ����j�WZ�)f��<�e0X�v��?M�0��@�L�Л�U���(8�NT(�Z���T�e�u�����~�L��_�Q�/V~��� �gkjk��A��&��*�c8�th�J����k��<i���73$�\[N���qqo���kZ&y}�!�"��A��t�- ����/fh[o5��9��_Eb�	���X��N�!mw����E᠋x��;��Eߜ�O�iha1���W��}Ti�I�1�m���j�J���bB� �z5�huw`ѶϘ��V0��E�Uھ�W����2	�s�@l��Ʈ�v����N�=��Za���+P�a�3Qê����~&O8��S�I�Pl���4�8BǶs9�
��:�f��b�馪� ҆ݑ ��	}zBX�����~�����5�]�;؀E^V�Ÿ�,}�%�t%GC?'���BZ���n�^DD$;����H��`^�\c���ڃ��gˢ� �O}N`��.H7�Q���Pl�6@������,�F�q���dES>����⌚N��0t����oP�hL�{(g�����L�Gmg�"b�v���WWW���`%�o��q�×�GD,�!��B�<�!�k��O��}}r9yy6$h�Hj���>ͭR�_1��x�e�i�����%XM�{�5�gz�-��W�zIV�ѓߠ 	*Ӕ�VD�o�^�Q	ڏ���(��54|����Z������@�^����F�����v3�,Q���=
�.Z��={V6¶
�_�$�cF(|߷���t����t�vQ�b w\���istPp�՝��=999�n��x���
�nA�������u�H����К��O+Դ-��C���n�AY^�8�״	x����!_\_ ' C�m�}�g_ҹ}�z��d!U���Zn���^��[˕���!�Or(�
���b0b��k4d�Β�>X*"n#ו�V�7
1��YA?�ѐ�-lp<�AZek=7��ߖ,�Q��(�"1٠��Y�<v)�/5���� �͡h����{_������^�,m�9�tb����[)��[�"�R������Ό ����~��nn�@>��� �	�cCb�f���!x3=����1�����p[��:��B��>m%%o]ϊ`�� ��X�=R�h�������� �:X���$�E*J .�.��x/�Zu�t�#!&�|�Pt�aoЖ�\8�]�@�>@9�,�[��8���sh5��V��tr�JZ�I<܍t�RS�C!+%��Z�B�a����_NҺM_{�q'5�+���(	"OL�$�>M� �M� %��A��PfD��2�����(����sK
ͳ��\�QS���G۟}�S
��ǋ�􈣥G]LBB5?f�PV���p[!�U�F�֢_��q|m�!��$m�A&p��iN�m{���0СZv�}���5���2�XLF��ZB�ދ���nF��M��?$���M�Du�Š�����P~�����Id�fmT~�2F[P\��7w���@�%��E������ȉR����u)-�@�����_h�7$9+�0A������`��x�A����`�bQhW+��8<�;&TU\yuB:��b�t�f�uz��N��Ih˰$�h�f�Ä�Ā��g������L�C������;�U
�����ܭ�H���1�9��}�EX�EK�%�/ ���ښ�o�Z*��ּ �2B�g��(�� 5��hn[��)��AVD�|�Am�9`a�]�4G@�U8��cͥ���	���D����i\����W+^��*ⶀ�dorX�AK�:}��v�f�*�ס8@Y;DOu�f �2M�D$�E���R���@_���V��[( �2�1��ͩ8t2�*��3��CGN�qb�V@��K~�*qe@����HuF��XNP3Ρ����((X+�L��` <���tP�@�P �4�62��q�)'4I$R�P���}��䙲*���RrmIV�{�FB�-W�W�?�o\oV�C��
_�K��Ÿ���o���x+E��r�7�*x�'Atc��s(M�4�����n{]7���5UKg(|t�Q�_�q��t�g�+���ڈC�l�W;�e�}G^�ԼB6-������݆	\#�JcQ� ,b�A�zL2g�1ڨ5�O(���$Z�M�f�}�
�6Z+v�/I1h�\ޭ d���@?����˦�«߀6����=��/�c/ɐS��t��N/�A7�6Kbo�voĮ`���6�JKK��X�^HHIm�%"�/��@vz�{�!�xy?΢S^��Fݕ�U��pq`�@��k�ɏ�K+�qژd���8h�(?��n���R�5O�VA�_V���%M�'��u�����k���9\��r�r��c��=z�h���
 �ZPc'DW Ovz
p��'�����D ��и5��q�_�i��9�F�bP$���ï#@��o ��2e'YMO�������#�)�
�s�h���*I�|0\LMt�h_($)�����n;�.�����?V`��j(�΃�;%N� i%������� ҭ�mG�����ǽk����H���nAU՞!�2�]�-ԴDR��Faa�7<0o�þu�x��Y�R����[�c�A�ʼ��H8h��T�?����˩�0n�N�1��j�(!�ۉ���C�=E9�>��^������S�&T�A�7c���v�I��J����hh��G5
'jk���P�ǕcT2�
�#�t��Z{,��5��nՅ 9^��St�����;�ɫ�?�����jS�� lhՈH�( ˶l�XD�.(�e�n}�("�0��*�P���(2D$�a�BD���s��<���W%7��s��|�x�s�vOll�B�j�{Fz':��?��<��d�;�n���444b�+�%����S�4��I������#��K��b� 	���ÿ�1V��ד����fRՃrL�z�#͡�Z����?�o�M��!���%��q���!;���5���[+�kF���H�讋�6k�� �ʡ�Y��<����Zz�^=��	n4���2����S/�}������ݙ<�@����O��.�C��8@���'�b�) �Z�L����㣦2kz���JR�*u����c��7�V�d�d�$�*\I�P�Ɲ;���5Zx�~_���w58�¬1R5�*�Aro ���bV�*���Z�K1
p\o��U�g�����X y·zRC �Z�П;0��%onV���V������'TH'	� ܲsR'�i�8O��¾M���P����<���6~&���j���#GV����r�V�\@r670��X3��U�{{F��]'�q�npE&%W9���Em���G�n.6@2ʉ߁QTOp%��A�HQ'�3�º/b&yi��F1Z�8�c���}O��l羾��Й$����\>����B�J{�y��م�$����>m�9p�߷5Ҁ����#߷Ot�2J�J­�֨��"B��B�`���_�%|#��d��r��z�w����њ�α��X9ڴ�{`�J�vrF�w��S�]C̽�+�8���[$���߹�I�L��I����>{oi�iIf,J񕖝�m��]�ï�YkH�Y��N^ ���d� )/|�/�R�dX��St,Z�`�ĭ-i}�@���N{r��SʟlXЖn�����,� d8�/�������+���2WB�G���ca�W���U���lv��T\�� �	0U$����F��1{NG$��s���4H�3\m���XQ�v�n����$��~�2ؿ��<���`!g%�SH6DtY'�7sETɅ ?%��1ɴ	���F�1��������?|�E�䐇Ė>���b�j�m�qP�+�+	�&������qݑi��,�ͽ���
P'��Ha��w�f�;;��<<�� $�Yӵ �f�3ݳ��.{��o��E鶧�Ѝ�+�����9&�p����~�,�ـY�G֬��qf)��xtZ}>2-a���@�f+G ��͜�\b ُb��������+:F��j�p.���� 6�Nn�솵��O^��e�6�����J�
�H���w� �RsK hY�����>,e!���f��;��Vlc�:�n=�
R]�!�[H��N�Ž���J�қ�-j�$<�:����VO���S�;����E{ƒ ��Y�F�ϥY��L�z{�!�F ��S�o���=��B�!������E�����б�F�r|F�pV}�gs/d+ʊl���C��M�ʳ
	�,��@�Y�Vг-P�GCL�!�~~�c����L�)̤!�B����!� �j(d����?��-|]���1���7���+ϚnlM(��̉CmC�;:w�e/��~Mׁ0�ۮ�/unq�\����a9��6)Oh;r�H^��/��dρ�&��c��q	G�/�
-o�A��(b�'�����p�"�N1�J��nԠ]����!y��&,�z�R�Hl�&���V�<1Lx%y����Pk��ZrL��wb�oz��c8�ϊ	�>ޗ�!mF���Ml��`7���'B8����lvf݈�{��Iq/`l[k�cNH{f��u��_�'�8 �;�Ly��D{�\���9Ґ�e塭5ڞF�<2A.����7�Ԡ��3-i$��[¿�	��YV�/���@������A������ui��ّ;��g��D�Mƍ����\�����c�Ϲ��߶�P�?y��˴�.�1S��<��F���5���W�^mV̚Odw����2-Q��p�Ih^Bd^�$���$�~�"�Y)5ѓ:t�h1�*��H�p�mQ�n�}@�v&�Չ�jtd>&�,!3�z�apH@P�F$i'6�e�@�GogH����I�;�`qz��y=]2b��fa݁��~�$����n��P`V����J:j��Ǵ�nbP��|�����L�@C}�e�DV��קf�k�!"�y2�՛K�u��0^/a0T%y�7��:@fu^w�
�.�Y�������Nu)�>B�;l�V��t<�B�K�3!��/II� �].�8�.�FA���N+��&�#�\I�~�"���H9G��h���#�/�qu�fu�ܨ�#/�kz8:U���)�L"��"�-��=M14G��e�p���CU���Uu~�H�-�Ԭ���r�	GEM#���#8G}� �k�����'/�|1s���h��r��*�$��	��(���%|q3�9V�{�x��{"��ɔ6�}����<4��T�F��B�hK�������ȏ�Ν���Auܷ����j��ޓm!�$=���^�'{�3�-��;q���G�p��W������npϢ���Vn�m+�B���hiS$ϛT�v(���R��!M}iT��*�8�-��IC���X�[��W��J�f`�9����ʊ�BҍfQ#�0�K��2[KK�4�)m�੯'�s��3�ι�����1n���ҩ�sK�,��X�}n�؍|��x�<�.�g�"ZD�p��А�Վ�ېJȧ������h���c��e� ��{ ��*A�9��/?�����`-.W�
#�}
s\�m������1�36�(��	��=����w�3�L��)����<?��d�bʙtY
��!�UC:����f�L�̙��0J�U<��V$㝈Ŭ�;���%H��@�;#B=+����+U�&��%�{Z��n`d,�R/��g��	b�=hҽ��ݰ��тS�������(�I�R=�6_�MJ61����Ȱvp�z�l@l;~ �WX�Y�'����`���տ}�puu��a��<���ei)�G��P��,������!��G�PDd)��[�r\b�>j�)�H(]9���.��֚�_J>og���]�*=����s�vl�+t�[E����ܛT���K��4@���I�PJ��|�g��#��Bm�����b����+��zޭ%k�WY{@4���1t�Ԡ����Xxh��|CC騄���!��<A6/u�ȑVAѳ]���b��sRj!�C��Y��nɀ�`�hY�Li����Y�$p�<��5B�_HO� Z���?����u����ai���Ą��� �EzRgv	�5k����|0�E��������t�8�0v�!6T{�uv�x���~T_(��v����`�VB�|�3��j�aO���� �]0 %_!*0-��D��c7$���
�B��, <߂ceRb�3Tv,�J�����.ZE0-����"��1����#��W!��]���~���<�R��*�LA�i�_��-=.Eۂ:��R����h}�}td;����d�I��>��	������[��Y�g�b��k1)m*���i�<ǭ�'*0��b���Tz��&��Y"m�k�d��uMl?N�J?�b�����{�r��Ԯ�\��������Vm+S��[V:h/���Hl�C�Dt�
+��K��Il����N �6��$��h
x��=1�*d��/鲣�P=#�%���4ߴ'��%2����V�Ỏ�ДY"���>�����"��v���LJ�\;	2�!_�j���+��s���9�Im�L?l�Z��I7o��?~�U4z�.SCz�r�\<kzd���#�A�,�F��9���JMM�����t����o3w��X#i���Ga[�?zZ�V̾�n{��s��DD1��K��@ ��<q~�������V_�v��^㤰���fy��k����u�������'֕$���c�ͷ���g�
\��ܟ����^BL�$�.ax2{)^��#7'��-hr�ߵk�J��|�z�!b=�ʊ������D�A�`�z -��Y��\$k�ų�~��Lw�$�"f:�4�U/ͿO��JDW�e���'L{��$$�,==i��jǩ~� �a�2F�m�_����=-�y��|��Ӌ��o�G
U����P�C@จ��o<����U��[y�U|,N`D&k�Q�е�̢�&��̓ˡ�����{ɭkZ� ��w��%���P�S�l��h�����\|�����1J`��C�o���޽��^]�����LAC�&$�+�7�����;��԰�As"���=3�"��U�"�/"�"3E�"S���B�A���Z4��KT"cPź�_#�Z�Y���C�p�L�wӽ#S@K�Τ��N��� W�P[7���!�������Z��C_텍�g�J �*�Ny"wЊ~��>&p�b��M��[y��Y���S�Y=o�zk?�3��������j)��ﳤ{�T�v<|��Hs#�A��#=��cd�Kn{���wĢ����aYkc����*)3;az��3��N�&��V���3�g�(���R�DY�<�j�J��ˤ���̍�F�ƭ0,S���X���A[����Y�m�v����ۧꨓbm2mW^s~��0�ۄ���`C��|���9�}��'�})�|`�P�!)��v��,8[�s�W���\�QF9�P��Bx
�!�^�.�XI�K�����q���I`�����_@5�L/R�ۭP�4���--���CJyE��>Q����#G']�:ZEc}���8���1�;�p�6�'r�JP ��$��:4�y�r�1���fLS}}`/E1�A���AA^?:: �y���^��a`����ɞ2�w����h�؀78յs�����팘^��2n�^��$i{��^A�������A�qY�]���6L"|��K���G�OS���lے��#5XNl5��޽{�b�x��&�Ǝ���w���]�X�_��R�D��$=��g���"��$r�[Q���z�K�jMK��	e��q�Y2�9o�<{O<��"�=K1�H�����E�e"?���[����٤�S%
�d:�S1�Od^�x�a(��U�ۖNOYEf��!jc����Rm�"d�1�o*�@^�uH�~��i�<�j���7�m������39f��Q7B���9�<F�5ՙ?S��2N�O�b�5onwf�C�,QoݫH�!�0�l��i�ɣ�}ן�z����lTd� �?ծ��D�������υҷ|S���}Ə !}�p��D���vi@oS�~��)� (c�~T"b�?�	�7mڴb���bF��e=P�bW~�e�zm�����Bz��(l�@��l,���H��l608S`�V�����4�D�7�0����C�d����K�����C;)��%;�����ߥ����\.���*��u&�J$�԰��'����_0��sK�~;Cq��f�?Կ�������23Ť�ِ���]�ic����󕞹@d�%�RO$���3������=-��'�b����j˨�(������"|^����|���-���y�砯<+�:&�j�*��������������3^M�'�If!ũ�~�!=��KC�$��xUm�VL���!A������b0i´؃���[B(%� ~�Xob#�Q�u��̩���,"fB�se��4������&�
c�^���=딏����W'�_�d�P�7�evD��N��<����EGH��Ԏ�~O��i�rAt��'�&��x`~c�{t7~��z�3��~�|T�.k?D��7��n�r����g�crp�!H����-�I-�[ๆ_����7��z? �\t��xlHu�h65!K��<E�_yz�#�^�ٴ����"�P'�h��,-U�>��a�~A`βr�txl�	�~�4@����F/���$��]�Ł�ԡqb�������({"� ?<g4�S|���¼A偅�����qu7�N���S�:�Ȝ���)�х�~�X巷���sfe�^�c���?���l�����˭D7l/�쎚�d�_.��ߩ�s}sV0���tj�P�)jz-��������~ ��.��A�]�R]z�\g��+] ���p�<��|
B��]��.��s����SdG���'U��r~���"ks�%����A/Ÿ����<H��]��4}��:������
��5��8CZ���3p�r�?���tK~f���EO�o���Ȫ��-��}�%���ƻ��ԺsC<����Θ��'����I+o��1�qo�2��"�.�ųH�[<��	,�8N��K����!ĉ�֏����v�8��(�����#Ky`d�����u�*ю�������s�q�� XI����p=�&f1�cG�(��*�5�e�����r�ܒy@oUѦ�#�Q�>����BQM�����FԶ,˺3��N_�O/ ֔���ݑY,-)\�hJ��rj��=,�'�ߎ�$`Y���o�_�>߬D�:��*$a+�?�E����$_.�1�v-`0�V�����Tk���xv|H�`N�n�\�^̑�s����%��w!tB]5�������f��l@�b~'����ru��ˆ�v���2���C����3Z���ѥ�u��>��է�r '����-�b�)]&��`��:�xS�.l8�y�T��w#��1����g����ͅ)gMA3Q�a�fQ�{�P����zg��6���� ��l� ����h1�N8pqp�����a�杻v=�c�.���a#��w˻�SR���ּNM� 6�d��"�}ҟ[;�-�V%<�<?HsL�5�0�?tǺӝw \(������G�r	#���ϟFcŨZ���e�-U=C�H��Nk��.�e�7u�̳C+�����u��������5�=���L�Ѻ�X���#G��	A�۠�xBU]����1�>M��<�Q(z��$"ڱ1|X8Zo���]��ps�MT����9z\�v-d9�А�N1h�R�	�P����<J���q�=�
�N����b{�%��!ێHKg��+��͛���f%������i|
R7{�����aZ���Di>W]�9�:��M��P�����Ԅ�ށ杮KF�]f�7�B��5�,��'ϋ��ģ\Jއt�L:��y�f�\�nQnn��2b�|����B��J4�c��p??�V��o/���hJ<�ߨ��wl d�nD3zb��x�֭[Co,�4���K44?Ɂ��0�D�{������S�\�ʯ��QA\�YHrU�[OX����~"�p��f���3��v_UoMT���� ��l���f55�Z��(��l�cJ��g�）�H����Kb ��*�}�������-|]�KI�&k�^�P(��*�������mC�SW(U���k� ���7�0���/@�KDv?u_ ��@�PtM��f��a�Y.Z�(��k/P�����Ϡ��p�9��I�9bJ��|�Z���l��	��4���scM�RH%��$�)0X�0�㲗=�gG�BG顤U�ӝ��h��N�%F�B�)��j�n���;f������`�ɬ�j:�;ml�w��򩻵��
󚆫+**4�lb�����T c�a#�A}7�r�0�͖�C.�Yw�ޭI,N�w����o���^|���?�V��HuA�iUY�'�6iū$���(��Y��Ь[]�:�ԋ�0�5�k�P����C�	�_��T	ވ��S��o�����Ϗ��8���2����tde���@WU��1-�cs�D��}��z�Λߡ�)9�%�71Z����"!�Y"��d/�V��]Ҕs��!w�<��_�1n�����e �\!m��QȨ��[!��	�	�Ro�>|�1�V�r|���ǌ�5����Ϛ�dee�!nQ8�Qq��0&S�-��e��D��n�52����l)��/��b��2V�l��P�M�C�����9[?/��X,^�Ou�c�{ޔވm<�޶��C�p%v��Jݞ�E�n����xb�VH���'o��tp��@���ng�|���.���n�أ�7��x ��x�-�����k���UN:Q����� ��7���R[I�1@Ԗ=��e�!�Re\�]
|s�ʃz��j��ё��ųS��4�R3�:�[-�(t�Z$v �����k�.Z�J���%��.��j���W�L2��Ԥ97n�:@�$�����Z�f��`qQ>����
�a<�iI��.�����~T�(y��� ��*��߹<����㍘��/�Txм掠�� "�)ڤ�x8���1B5�Zw���ˠ��Q���r����h�S�'v�$Y��W��\PP0��;x����2��E5����A}|����@�� ������u�qn��\<�)�a?Gy��c �t]��Q�D�l�e�-�~��rW�NޡE+�Ju���`�;����!�Y5��t;ā)XUB��Gr���%pÉ�#� �X�YoHߡ��S<��')�e4Y諌�������CS��duc,mx�;j�9r�#)�%���B��eD~u6]<�ooB[yV?A[�(s����� ��o�!�;v@8����`yRrl�;e�E�Z�8�f���P�C"}h�#;D��s?Fk,Y����w+66v�*��a��@CC�	�Ԡ/1-���UU�%�F\8�*�hS+��i�K�����������69ʫ�
<��A ߉2���6m�8��=���9�bJ3��&��xъ��@���Esk^"��Q9g3X�{rݖ0�ȘU�u�I�V̘6�(W�6�S��?-�٤ &����e�#2�#;��u��.ʮ U끠�)7c��/����}����������4����Ё�b���a�a'�vݘ��g���aa�(���tv�8�(�BT����0��D�w&������mp�����}ׄ�����P狁n��6V�ǜ�#�m�h��1���C���:㍑����x"����H�5�ږTP�9�ʸiݙ����#h <R)cz5a�����{b��.Yz�oò����z:F�LJ��7�Y�q'1�5h/�)rI�%����ץE�B��hMݩ��i<��6w��Yu$?m�����T���ߤF�3]d�D'��{���>��EM�P>Z��q!T�_�ñ�̊�<QT�*S�1�@���F��w� �o��2e�y���:
f6��ai5C���՞)X����H%H��|��3�mb|,ެ$	�\��4�A<���2�ʠ��Ϟ=���VhİO�=��w@L��?�+�m��D��,������H"��ug�I�5�J�v����CG�U�P���V��u��(k㯮!�Ɖ~�r�?!�Ӥ�m�b�����]�?ae��2�)��C��|��`b��xOHּp��N]�z�Çjݒ��3�@+�n�p���;;ZP�Wz��z�ׂ�O�d��\��(u?�˛)u�����첔�
X�������}f�
��v�.D�2B�_8CE"Qfy�'�Њ�ֶ�=򠪫�j!k�ۍ=�q{�(�*]%�(6ԡ=���{�c}���L�$�����&��ai��Ό���(�e}��zȝ��A��D}la
B�A��[A�%]FK��aЛ�i|�?�U�W�u�þc����A��:uDx'�cj�+�A�tY$�V��CFffx0XjՖr\�7�"䷌��%S��3#�#P�#�m����mN2�Tϸ�f(����g�m���L�1/SU+z{)*�7;]q]]�6hmI%���vG*T/���ˡ�K���H�+)#mV�5=m��Ѩ�H��nUi�l��ٌ���P�:֚y���IrCÄ�v�Z�SMAC2��Ua'�K2LJ, �ǉ�_CI�ɯ�z��:��:TmQ���J��BE�ж���iGQs��mݛ�Q��դm���(k�#��{��ŭ������j-�c�T뷸�U�_dRRK�{3�u�/�鮯)���6��ߒ�sH�[�x�ྜྷ��맮Xg�@����o��g+!�y���uG-
�>�!�1�K�%j��e�"�k o�'Q3��{��y��G�?"�����oZ�v�
��Ɛ�� ��JMK��^�7o^�9PzV�[���?\9,�����*����L?���פa��gcT(��g�V�׼�C�����.Doo��u��ug,]G�z�0��Z#��Ep��'��3aX���`���i�P!:�BF���:��(��jpʺs���̀��F1UH,�ynn�~֕	ԁ��Pw��*h�Y��16�H$�2z��R��c��S]N>���CI���^�q�����^�nC4G�lw-���1}���t�=���s�"�,9C���� ��5��<]6�UFk��,=iz�3�.���5ϵ+��
�U�6H)B���,�0�� ��EwI�Y�toB�9!}P�D�Q���U�އ�q܁)}E���RKgM���v`�؁s(B�}��W�E��*x����*�V�� ��1c��D��Cew^�;v��c$+ӓp]��E�x�4$��H���t+E���UZ�����"��ٿ%�w��N>Za��5 �H!����tz�II)pQ��΂�������U�?|-��Vs�0�Г�k_�X׆ҥ��:P��eR�y�h��Ћ�\�������Oz�|���?O��YJO�*�e����C+��r���<y�{EdO��a߲]�w����9)ݪ�� Wa�� ڒ�����3h��(���w��{�m���E۷2�ēP�v|�%�9����#Z}p�B(������7��f6m�QәF��R���N��N]�쨾lV�	~�r�r���T�0�������@t>��hŇ)7fݾ=<b
B��;i/݋��6�1�ڕ���߇Xw�-@c0���aF�x�V�����NO.굄RJͼf������Jn�����q����W�?^���jn}�GfHp�������@��wіn̬`�}���C������s��U��S�;�l��JW�j�i;�m�w/��55�Ӳ�2OpF�kb+g���4�6�-�V[�G��3�q���ÉG�Y��Y7��8�[�cI�>��H�v5��ܜ��
�<n��fp�ԝ�98�8ȝ݀O���d�O<>}�I�~�]���|�II(�k��6/7�?9�����MvM���@��}~���p�O���q�Ol7�%� �^;��S@CT^�:Q�
��7�\O�޷a4	�]GP~σ�ל.kP��W�~������Kb�"���6::ڳ<�=i��P���[D��j̄@��L��i�$7�Κx����V�,J;U�Z�(��!PVD	�w7M܂��xt
�ߘ�4X�6"�S_�})�b��5��J��J �*���b�R����)����T��ž�|�W�u��R��Z8k��H��WU���&MT���C+,����n��j�G/l4_�5��J�����2�	Ɣ�ָ��t�7��G �����ne려Zĸ~���!�L�F����������e&%��Etls5-(蕁��L�mڦM�R��',E��5�0Z��ɩ�?�=�u��2n �j���A]��E!��G�]~Yv~�������~wwwC�Gmj�T(�`���dH�b-
��ֈ��)�EB��}n�y�[��Z�h/�;��͘Z�6�;��:�+z
��RfۮP�P�_�^,c�A�
x��*�����xA�k,) ��E���>�m��e��S�Om�82V�����������F���0��{�w� -'l��ԉŅ��?�.%-�T�{�{S���GވBԍ��Z<��LJ�*�>vuJr)�x�/���ݻ`V���(I������|
��6wdk$I�zVƛ㬯"'gPvo	�N>��:�xiii�A�>A��:QX��X�h���d�4`Q���EY<&ވ#�})��0�L��؉�_�Q5�o3�IwI�h��͘�(à{P�z�uT2�Y/^С�I/�c�;�w�^��G��T_(K�%��{c��?�0��_W�^(~��A�����%�q*G��E�ˁ/���52af�C��9�����e؟"|�Ỿ�YؑJ#|,8W������'��ms-x�8$��r귁h�/Y����P����S��F �y$��OEn/�VV[����#��IC`����d&ɇf@9��H�~��h�öQۮ���΁R5�]b�3%��ۦ�c�ju^��Tߣ����]s}r��V|�䖋�:R��1�ut�9Ʀ���(uG<܋�m��th��:^@�:��b����~S���U>�܂c�s��Ռ0&n#��*�-�15(q������� Ӓ^<��U�I�)z�/�9�x�}rCSS�zEg�+CBD�ƩM�]�z5�ڵ`���u�
�o��Yˀ�j'�"�=ɳh�_{Y�G&�Ώg�v�♧]5v?i����q����[�Qs�{��ʶ��E������;ߧr����"�Î{�ά������_fݢ3���_�j�����]�q`��}Ng��+�/�R��<���ƒ{_��h5��j���8}.d5�(P�u����r��8冎k��na�0���s@��`;F%�ŅI[�4�eH/�����s�D�75@C�\$�3Z��T�<r��0,��Ra�fq�}�X,�d�:��6�U��|Ap�1� ڠi���!M�x�0�o��#�¨�.��}����5h��:F�-�{13��d�/$��By%�/�P�rL���E��;�,; ,B_��s��2�.0�	��a�	M�q��Dq�z(D�=a�Q�60)���&��]�Z����=���]��Dw���}\#��������+�j}C�?ѳX����C����������u/�{��:t@hܜ��;0��Q�^���*��W=��贺1>J�9�Ժ��0�Q<Hd���3�OŻ}�U!99�<����('JU���{|||���e!���a����J�)/x:mI��I�z\���9ja�� O�P����gόc-��2�QV���o�)�]?�݉�V=���M�5 1u���L	#�Ip�$�� �8� k��O7����ar���@��OBnS�#��8W5-�ka���a��X��T\�,���l�blw3�0���)��:|��,����]�z}S(��ߢ�5Ƽq�[�9������(�e}����)�g������}QSq���{n9��ȸ��(�@ʯ���"��|�C�71�V	�`���7�?�m�\^��S$��5|b-�Fޜ�z��3�������| ����WGa��d�7v��"�,ժ����Ng�fv@�x��%�6݌����
v��e�C!~Ѡ�	e�# �Bk�9'��D��vI�����
*rp����`d��7Gu�P�d���=euHS\���N:�b��g�61�LJ��X�"�"d�)!YK�>.���Q8۬]̶Ԯ�T7����K�+��)��0�C(��r����EЧ���6S+0B�N�Ѧ��K� k2dl���������*���'��a�Wa�/W�}���R]���u`�/F� )��O�r^8����gڢ����f5��e(@B'�x	v(�Λڟ����ݵ6�*V_�?8x���T0���yi�����o��
��y���y��+;��G/�v�:�L��k�Ǣ��������{ø�8��\�����@�����k`������'������*�Er�w���՗K	 S����sZ��E�rsv�6B��!�"��C+55�(�|�L�(���o���-��w��r%^��2�F��_��4�K��@+�c8r���|z�]_-ڴH����Xͳ8�_�o"�����Q��20�7��g��w��2�F�SN��0������nb�T��'Х����a�y�j��V�u['�r%�\n��P>��d�� '����#L��Cv��4ۣP��Po퀝�����u8��-���Ŀ0'��47��y�r(��6�z׮�-�R��j�dqMP�L��t���*�=˞�(��t����1f%���샵�Vk �S�h��eee/C�����VP�Xa
0D��8����vΐ��c�o��S��u�j��r�@�?>�T��O����#����7X���ao9螺?�V�J�DO�c(�7��W�S�̀�ĉ٦N�F��ns]����6��d�Yǂa��������%��'����+���R�D����$G$�WX=��wW���)P'!��N�/�}؀J�����E ƒ).�ʆLo�&�.�
���}�ԗŹ�/�7�=�OL/W���R�5'�������.�u)U�� �zv��17�/���ۦSǓh�?Kr3!�籟��~���wa��"�d�Z��6�7��}�;�1*������|3[���ޖ��S�'�LA�����9Cl������T���v�L�)n���#��v��O�:]f
���6�E�}�>lt�b���y^%B̒����\�e#��c�Ae��������\]T�H�_�����[��ݻs֮I��ܦQyMŻѯ�p�r��}�	GJO�1j�窤��
��"�����������+���̢��6aڌ�+�J��>�h�H��ԗWoڴis��3��~>P��0C(.�O��F܍Rbr����%ɚ>��غ��!�[kS�8��%-��u,V����X�.����8�)8�ywC�e�e�� �GP.��;T_ҵ��-�K���6�O�M��S��c�p ��|��q]��� D���}��9�]R~!�e]�͚������m�q��&[�?:��� PK   SH�XN�v4	� m� /   images/91e5cd07-2a88-4b0d-9128-72e2f992e16c.png�{eT]�����ˠ��Kp	 �Cpw$�%H ��'��Kpwܝ�y��_{���9s���vUݺ%OU߉��*��F�  0d4  j  � ��B:��Bt�R��`�H�oT=w �P����S�^�����t���6s�X�Y�Z�[8;�譅�(ʼ��u�����.q6�n5&��h��H��tҠ��_���o_���ݰj�9�j`@LT_�Z��d���BX��%����T�^�O?�ڻ������;�^�t��#{{Thm�+��j���J;�?��G,d���)���'eH8����%cG��q,%5'��O�N-J��dj, 4��v8?Y#�0Ӎ��?�`.�V��z1�O�������{W�8�^����ap4/~b^���P��^���}��@��-:P��:{1��ΑW LQQ���Z?���U>�Z���N�1C�]ɅS7�HM�3���?�Y0��sZ�ۅ'� ���%,҄nl!���wD���`G�b+��O�~������)����,�J��z Rɻ$�-�TR�*Q8=g��?�Ѵ�Y iEH$#'Iz�oY����+�a8=��b0ҟ�B�T��}��;5ʻ�;$"�;W�P��$⛩�4�_g�,�� (7?�Ɣx0@b��awr��`��1hdb�Ծr����Cq�Ӿή*�Ä�݋�q����LR��\�v�Bo�`�z�̐��I,���F�4�!�����!�
@�p3O�ij���0.����ZeE"�X�%<|)�ؤ!�`3�2����a�ƈH?��¸�$�� ؈�H�QGjC�T�ژ�B�`̄y�#����vm&��"��[B��IL����g"����RhY-��C	�
�I�H�VAt2�w
�Z5����얜����e���!V�?���>4���>*$��H՚�n�	�RBx3N�K�#�u��_�u�a$����8�d D��1�J3 7I�*E�ưdB�������ʠ�DJ�~7�S���yj�d,�8#V��K����������,�cʪ�c��C�������b��Z�8]| d���f���g���sj�=�� ��x��!�&1�r�Ӕ�`�co����#��&�Q2G	��~��^klQ�0>�s�5d g�B=�d�H?�JsVP���/�ama��&��?X5]�(b�Y���ӣ@��w���'�.�7igi੅�)0��VK��E�i*W]�Tu;=�,����?��7q.N�;�.��ڴ�[P�B�6��[T����*.E��ہ-��'_sI4�Ҡ����:���=8R���	*�+��t�}�k���7b����{��>҉"�T>CG����WV�Z�����Qʈ��^�	�?��9�̫P/H�"��w�Z�S�;WT�x�6��:��I�R��E���� W�}�}�{�*К�ì{6\m��%k5'u�A�lK������l�	u��4�x�J�r��
e"
��ו�+)�3�+�֔�OhԠЏǻ��qF
.�^�TȦ<�dJj�_y�8=r�v��g�E���0�ۆSkJY���{��u_�#��H
߾��92��8���� R�b~�4u1p�iF����".pP��j���{�<���ٿ��Pu��,���t�ڰ)կ����ݵ̷��xv�լ)���;f��h�N�y��?���=E,��&&���;�"j2y�0R�H���)d�����m ؉����3�.� �U���ցm�l'�2y�1����&T�70vႝU_�X*�X��ˁܟ룽�����<׋y(a�Bᇇ��|�է�/�Vē�'�)�o��@i�_Gx�����I�UeO�Tl��	j��#��Q�TӃkw���G�C�#�X�ƛ9����2 j����J�xQ�eC� H�X�f����t��tPԯw�A�n�r�7}���R��uNOǈŜ.�{����U��	��z��잤�a;��ب	��2;�<�U���[�0�6CZ�zP ��$�;�k���1�����-��&}��ܢ�}2Bsh�쫠R㥭=�?��65$꧲
�Ɏ"|��b��{����|���M��^�$�0 q�$"��Yo�Mp�+�ڊ2�#⫩�+�>�����J��t+��)�W<!��K<^�>�ې���YO=����Q�%�rpb�Q\G�vË}il�
;͕`N����Ml���`Q�昷�;��O�S̯��O��R�>�}�Jwɑ��mq^���Z��o
~p�EI�DŢ7��M�������SI��C�2�YWT�N�I���#��
O�1 H4��\ԶP��@�^bG�A6~/h�N�K��'����"��Uo3�0��i�ZI9V~�9�(�<�Yk!fӁ�4B��e���%�jכ'>�4��?Hĉؓ��8�tˣw|�AbH*:�I��-FѴ�����M��.�����`�(S>��H���ϳ�� 3�m�j�=�r��.��fm9�B���!�+�nc�x��#�*����k�S�B�������ug�.U��?_�}$J���wB�`\��PL%���17���/���[�YS>n� 0^C2 hs��Vw���/l|���!��}#Vs�s�㐻W25��G���c��޷Y���LU��P�&�:����-|ԩX�z�Z��WM;W���*l��@;���Mc���x-s�������k�*��}��Y`}��� Mx3B�CU��_�:������N�%��WO^��b�*�z�oə�h�B�cNE��<���½׷N_�}�������ڑ�)^���L27oL��Bj�q��Ǒ�9��=(�}���s���=��D��	.<G����ׅ�!�8��t�v;ń2��Dc{C�-Q�g&#SN���Ō��_ -M
�㘑8]U����N�˳6���/E�`�G��f�eG�q���0C���g��2��JY�!>r�D�]
���~Ӷ�$x�H��C$c�pG%�]��� ��,��q���=5�f)a���1h*k^��G� >�s�bQ�E^��J����1�uYL�:�
���'��s�!�9q?j6\(�x}��c��"_�[C?i<=���)�v�e�Uhy�Q~�g��
]������F+9F�8�FƐ,�D��觬�B�.�1	�?O�y(�D��y�Y��"�P\��<�[s����c�U��ߙ�*Z?�H3R�C*Q�����-ȁ���*7�HN���^gA�또�s�����`U�D�mɩ�V�-����i
z�8G0�U�d��;�H���X�95��YE�*�y�Ħd�{|ej2}�� ��Nd��tw�"t�h7���"(�2�c�G��ɩMb�jj�t#a�G�����A&��!�Ԧ'�b�l(��E��4&2;��l�(>T靳�.N �+�F�����U�;��}�mv^�2�vd�Ϋ�%���N~���d��\��U���=�����3��]b^~?++�����3�1���8���
�i����d�H�K��Ѝgb���I �5���ҷ}+.�
&��!�25���Ք&Fa�7�0@�_����}�"Nl+�q���/��&qY���G�5�?(*�5fvD)TP�J�S�Ȉ��PW<R#>Y���W�l����<+V �BE����֜w��]�/؛.��ׂ��{�K�ޤ� EO8[+��Ӽ� �)+��4ro���T��`!��'��%�յ�::� cc�ٙ�M8��g��J�t-���k�ja]�~9:�k�W����t�+��$�]C�3��i�޹��F��=E5�Smi�?�ib�3����<ȯw|�����^�|�^D�7��[�]]j޻K	$Á�P��&(�MT��"�6r%O	�|ԯǳ'
�7-���;_���κ�9ME)zJ��������Zc�T�������7P�Lʀ�DyP	\�Hw2ny��S���J@��E(r�e��Wɾ�����s�R����E��36:duǩ�bĖ�*��~���i���}��;`''œ�§��Ξ���{�5���ɶ�%�Aj��K6��rባ����t��A�x��9��{�i�tCk���D�ٍ���a]��Q��_L3��|�wϥ��[Pp@�G�2
>�ʁE��F>�N�\Tzq�Ҋ� ���#`Ax��<)h��N`\���A�6���ċA���.	��-UȈ������ἐG=-�|xȤ��9�����-�q��[�?�~�!�v�;���;M����O-���Ѐ��3�HM=q�/{!c�� `���|�ү�*OK��0M�t���"*����_,�U/�������/�NM@�n��_g5�7Pi-,3�$�J��z�#r���H�#�'&l�ΰ��D�8U����2i,����V��{#8pB%���eq}�쉻�� k:PJ�Q�C\��𙦟�
���F�=cI��lv&�^��Ɍ��~�Նc���D��m����fWr�P�*�Ƅ�&�L�+��'U��¼�sB_�:`�ɯ	���S>���/Y��cG�vK�O� 8���>|Q~	�頳����p�� �.�k:	z	g �Wq��5r��k���?(�k���R����z�����=�bR3u�%H'v��~����]��'cd��;��֭��G,(y�����U������AVc�m��}�Y!�\�uL��P�b�;�Lyr��Q�"�T:u?��$`���^	�]T���WF�����1�[�����1����l<}<$�i�@2u����`��5��ù�p�\RII #��Xe��i\N���j�X�k?k�R���]���^�pa�x63 ��IYd��HI��&��!vy�o��֩����,�]1���K�}�������8����J���7����j�������u���+��u�$v	���F�eo����J��G+�9\��c��_*q��>����w
��S]f���٪|���(h8Q�D^�:������E�'�e �?�7�e	Pn���I*6�|s�W%�B4s����E<���Ĩp�S�w)��:��@5��솢���YPH2U$�&hh��;���k!tv|c���+�s�h�u��"�]+g��w�TQp��̔�=��k6�>ǡ�k,!�+TEWY �%�b�[/̀�������2&ȍX�*uY� �z-��K�h)6/Q��1���)��Kbldӡ6˟�@ַ��� /�IHۺP�gO��,���|���M�LQ;��7��� ��ޙ�-�x���o����V(Y���ܿ���S�)���i�D��}lY��*6���괷�Ľr���x����.��2S�]k<����G!�u:������AD�8S:"�Y��||�'��O���,$�Z�6C	��X�HD��)}!Hvʉ�5�@C�p��p{b�ň�H|�
��B�}AlJS»k/���^���_��#��}G]�&�6uN+�o~^��0��mQ���G%��[�ö�����r�~��C5�������ͪu��ֻ��%Ց�:�����J��UD}�06��=�[���EjɊ7O�]�F���?��u�-ř��k�V����s���I�<x)q�`"��{J����a.|%=:Ol34��+T
��zK��sN��<���2��g3��6�a��м��� �T�/��s���:}o�G�AE�cQ����o��i��i�`#���\�&W�=�h�/.��قIR@�Z���<�m�ݢ }����15�\�h&fk]�A�ۧ~'�ڑ�CKn[����H�x���� �Q�|�����S$�%�M���bgu~/�@*�3�&�rQZ���HL}�G.,>�g���栊LB�'%e�ԡ`+���X{�(�N�9"��U�~�3�W��?v���"wYz�dρ��w�BJ�̅_�&�7����k��pxMnй�9te^+����@��e��ȕ�o��M��\x|�iW�A�S�'���N-�B#Iq�+K���oY��WeL��OMD��\�<?�nu�>�)��y,�Τa�>w�t
:q��� ���6����!)���c���Q+�u%��p�-��̀��{��#]�p�iI���Ϋ�cR��b�6��ѩ��!��b���O+�b^��|ޭ�PP����*�B|�b��H�{>��}�S��.�Ć�^>O���m��`G1a��HĬy[�LAL�:��V��u% me��P��Tw)%AF�(,��`M 1��^�>�D���-ə��,]���ȩP�Y7���u���C�6�9��4B���>IƐE�v�;'H��2�.��+����j^���;cZ]�Łb�c�;�"��UT��G9������ij.T5�����'����j��k�98bu��o�"���ۮ��RLb@����Qv���,�$pCJ};x7�	6SN%�=�jw����$Z�h�t+��S�̇B/u�B�R�9��2��W9�t�t�.�TJx����)�6^�Q�;Z�i�%��͗e�m��1D��ߧ���ı���y	����#��px[I �� y������)$��4��8��-q�5�=fHz�z@�� �z;����#�ȫ�����jNF��K�I��7�)S�K�V��#���?�?�[����R>����g��9# g�'�~��_jZ;�V@1h�I7�?X��֧��H�Sr کh���*��"�Gb��\T
B���Pq����gek_��x�9�q���H<�iV^�~�_)�B�E�ANW�A�ːKU(N��Z�ﳂ�L
,�[5���P�Sr��N�Twʇ�[sq��D�λ��Ռ�0�����y^���Þ���4���T��U�h���w����>�{�[�c��W!@j�476�B��m�  �t�w�:�G�@B�&��TVXk�ͥr/��F�jВ�*�꩝>o�^�=PiN�cP�U^$�H��M����y������'8��ى��\k�W)�rw�~��+�(��K(ݸ�[��Ҫ��rYĄ�ԡ�&p��E���?άٝ�55��`�4=���O�hÞ���ϛ����лe?�K����/���M��,h�qB�w��5�oT��e�mq���8���k�j�`����BVU�3��e��e���C4�N8��&��p��+�Nd�Y���1��F�]�b��Q8g`}��lAx=,�AHng;Y>����G�Ga�5a��9jh֞�"���ڌ�bl�Es����rЮ�v�i��ٓ6�f��k�Qk�O҈���J'=�)8��Ԗ�.&n��y��&P�E����mc��]Z���x �~sc4���K�+0�LA�iz��Y��`|<���S^K��48�% �%���k,R�7&s�vx����)X
X��8��0D
�B�§���͈,ݒ��\P�T���R��I�`�U���i[`H"@=����S����}�q�=7�胵Fө�_�bo0kF�2���}u�ΘɁ~�G�B��6+��o�́sA�	.H� �|����"�k���;CRu�'�\��7G���
��#����Z�g~[��J�gyq6h��;�æ>�T}c��#�b��ێ�t��jɜ勷R�}���w��o��%s�`#�_�*J�u�>��us�P<[��#��X݄�Ћ��?��ce�G>vX&|A�1��-�!R��6,Pء��a8U�yY���ܡ�0ֈ�B3Ay��F�F�.ۣ�!����U�`��� 0`�W�Z� R�%ġ���孥8R�r���ͣ���E�����e�[4���؄~۰����/��]��f6�Nh��a���B<S�ݺ��z���w)�ЦgOսQ�!�hkN�ܨ����1�.���h�5���U�w4I-��7w}�(���sz����L�=!���r�Jf�å"xTe+^U�)�c��VcY��\O! �G�G�ZpDYY	��G�>�إD럜]�/���4�Z�\����UQa�i��_�F�B�Ǿ���$~FzXgв:����?�hU�J��#�`��YSk[�Ys���!�o�ꇻ��Џ{@T.)IU �|���g�~/��ij�Z@�iK� ��҅M��X�"M ��$&�o�O�1�8�*�܎��9% 1Fi��5Ź����qҹѻ �I���'��u<لc�- . �K��1I~Ħ.�A��?{�0�e�/��������qv�� H�4���v���Q��YHO�����`!Pe��'��st��^�^����GQ�����L�9Ro.��~�^�T@Ot���qrDـ�[6F&��j_ܜc�����P=l3�.���a���A�]E+�dN��޼�w�*�y��`�t�I"Y�v�W��Hhv��%�Ĳ�������-"�/ߡ{�A�b�%>Lfd�C|^f��]F��V�OB�/�U��,�:{L��k˂���W:@�7:���PÖ9�}�h<��@�6,u���F;M���[鈈d��H���m��Yq3��Ж jȣ�����+����ێ+�p�&�_�M[�(o����@G�=-�d�U�����*�pu����h��XV֦�4E���)���8ڮ���[.I�kdP��J��<�~b���k %x��{���v݅��\�~�(�\���;+�j�ix�;_�8o&���FK��� .3کB<�W�-һ�t� 6o�p1�i��޷�g��>�Fw�<\�>z�Z+G���s�|�|�e��Q�z�����{F�=����0m�B05�<�$���k��t�8����m[�%uY
l�$����J���� �u]B$i4Ch�E�1��]�_эCf�lcs�6�#\��%Ej�b���cQ��he(,�=��	�����1O37Ḻ��Yy|��wмE����V䤑�t��N0�a�J3?�������q8蓻֫��v\;��mE��0�H��?��-X{��
�����b�]@OB�����~���d�QLu�>X�f�����P���J~F��B-6��[��#]߳�1�oRl+|Y�o$�O�4��?
��J��������9�B�$���ʯ��V���F�Cɬh�4Pf�ϵ� ��D8�<�܄E{�;�k�]��e��d�A%`�=No�#ɉ��/6@#_��O]���4���(���F��Z0�Q��[ZwIss�d�O �)Ӿw��}bn1"�{vxwU��ŷ� (A_�i�#�m�������ӣ�ϲ'b���v�Iv�^N�ޘci@rM,�#n&s���6&w{'8a��{�Z*�/tAH%-q�,�h����϶�x���󚹯ߍ����#��=J��}Ύg³%F�zo'rC����U�d|$��V^�N����_��ZJ=��=�KlZ1�]r��?vtXc��OqYh1�e�:n��8�I���\Hi�.�{�9���[�NS<���w��o�ꮎ��Vۼ[3����R�?��\!�[8-bw�D����C���_���;huǼq������ro�C;F5��Ng���V�.|�"�D(\�ߧ�u���� H��y��1r<��Rֆ�]�֞��k�T�s�X�YRgU_ʡje�QX-� �4-#��u0J��+ɮC/(>�G�6a-4h˳F��o猙sՐ��ǒ9u�X'+&]�!��K%��~��},�m��"*�����c�·f*1u�ۭ�oo��}���yT��0"%�T�~�]��
��VTdÞ�(!@��k���1{�<��,��rY�5�=�
�V���l�U��"��E:����H���z绡1�w�N4ܵ��"�f��?���=�7�{6��*��D����VZI<U���i�s�W�3�c�ck���*�6]>�7!E?b�3ސ�d�lV���&x'�Y"�fQo��;W��۝�[<�em�y�&��/ʸ��'q��%���I���6���;������r�d����I3���^K��i^&�ԇ�o(�D�{Q~@e��W�*�	���)���D|����o��uQ�D.
��"��\ԁ��큮��[�1IA
���v�� :���<F�$�I�h���S�(��Y�M��Մ<��F,��\�g��ݒo��T.����w߄�LZ^U��5��c�w�
�DN�E��������A;Đ���>�����s��t��c�]q�>p�!aV�U`a0�b�v,�m:v�ٻ����軱W�������n���|�Z^�^���_�t�/���E��`��N��׎��؞_r��j���v�2?bŠ�D�u�� ѐDV�*a���!m�i���L�H��!�a3��/���ߓ�k�;(`W+ k���K��ETѿyv�����P��`���}+暘7<Ѩye�cS����P��*�$E���Cμ������\��ߙX��K+�*�0ȅ0C�s�V���'����J)f������4�՝~& J�جcILZ����6ɲ��H�Z�qD��4[�,�����Q:�iN�z�A�n�=�3e��4����m���?b=8�P�w���=Zl�E��$�ܮ��=��y=.5�/���6��b�J��#?ʀjN��ϳ�?���ęт3����ƨ��c�Ҳ��dL���HĜ��l�9Gۙs+*�8��a8Z��\8}�)�o�&`�r�R�	?n2�dWR�{�|Ya�Gr)|�Y>u��^��+YK�b,-���i�gRj<�{����]8���#�~�=� -��V�T�����8=3̴�.;��U:�;;�n�ii7%���Cд6�xʶ���m]���%T�]�����������b��":O�JV~/�^����=qЂн��	�Ш��olii;%�o�VVb��O���}n����=�Hcy��24ifap��B<���y��m��5/���v�5E�Egݾ�~��Ǔ���Ӣf�����{�&�Iz��N!T���0�|�${�Ϧ�w�`tŹ�pB�����4n�5��W�
C.2��r �s��Ɇ`0�JW�:rajo��E"���ÃR��B���=G���'Ku�ʋP�!s쳚8�J�P��>����Z{4�?6�[�{8V�����P�FVRTt�������y���5�ʲ�^1&HĞ���E}�-I�;,��A�S�%�P��U��v������M����d�D����%�	��k_�:{��TAoz�;�j�2 �����NB�w�O��lx2�Gd��1���b�A���H���]<Rw�>��#%|�����&O��D��|!f�ц���&gٸ扄f~�_�K�j������6Zy���:����̝Ij3�M�ojz|��b��6�P
�5c���a�}:�ڣ&��=qdiS��Ew'?�߅�>|�g"ͺ��n�Đ����U�� �ꚴk	�y���.]�^ň�������k��5t���(�ѝ2��4G�]�8xBa��2�7����<_Z|���ҍ1�;��u�n���}k��rU?�\�r�����ҍ�8<�/���7�7Z�M�G�$_3E�����N� A������hu���u�Z�K��̥fb�F�Qe��lk7�Y�7�[+!��u8����,�Wi�
i�h���Y~B�ţZ�F���N��@�}�/�o�րN-��aG��)��.ua���mRwҿ_��ϊSURrV�^�G�o�AB��~.���,J��vtk�ɛ�Ƿ�ht�ݦ�����ꕃ�c��6�H�M���\L ~�C�b����_C'C}ɤ:�W��TۺW�8�����A=k���#\��d�O�+9P��}�����?�{��D  I�iO0-�n/aX��׶~]>u�keo�H��B} ��ͳ4�Z��l��)@�5��.���I�M����
^,�q(��Bc���?�);�cOkQ1��x7��8W	5��/�&҅l�9|��:��?j�Ǧ[TpW"x��/}v��w)�����9��������썿Ͱ��qp�h���)!�="/ap�.5��GL��(�V�ty�O�{&�)J!ֆ��7=Y�V̧���MH���:��|A��0�+�vq�pM{O����Q�w��t	�]kr,��6�C��3c�ɑ˷�l=9e�㟔�}u�A��R�ѦZ�ˈ�[�_�#Օ��u��xw(�\,=::��m�h���)!qk<"�ی�/��.;�O�2ȏ���Y_�~U��~�}�ҹ j>�K��&�v���X�1�����w������g��J���������67�-�k��$)!y!c�?��7����9
�����]�����C�	j�����{
R/��]}�
�Y���K�^Y�y�5!��R)��A�*�����P�CH���g�T�,�&c��{t0L/D�r�(����<$Ѱ\���.��i���Ɋ��&!�8\��+�J��]9�˔�M "�=�a+����ԗ�u�h�I������8J~�����i3V���ÀM�F��S��FuA�L�x06Q����p	r�J�-�����Q0�%ay]��U`�?~arxPV��'V>َ��,p2FI$�y��dt]�T҂�	���7��� �!��P?Y�~Hs�	�.�{�ﰊ�wy��?#��3��Kc��|s#��#�����N~{.9���
.�H5X�|�f������ ���j0�#"�O������ó��vo_�q��p!�EB���ߓ�**j^�Pi+�Rffx1��%���I����n^#��}˝��O��"���!HܧI��r"��_����W���Q!�PRS�SW�Exxۯ�6�P���|�2��*�V�8ސ��-?�|_̶��o���OC�b�H�Љ�O��ϓ�5K��e#�#��;��!�7Ϫ��h�����zK��k.�&��*��U̾0�d��gƓ�[���%�j�7q��R�����Ó3����L� R?/Vh��kf���jL�Ui��L"�n��~�v!�j���0�.��e�����q��A�U�4@a���{R�E��D�۩���M!'�$�1�9N=����YVZej>��±��3�("�����+�����p~ޱ�r�`a�D6wV�e�D�IN6b�%��+*�������!+�9���n��
��$4pOfkr�n�m�Ld�zQ��$��q.b&�o�Mv���Ѩ��,�^�������q
�r�I��a���i������y�cG�ŏLt��˧���R��*�!b�G���	$�کO�^�u�1��Q��8Zݫ*F�z�Gp5��C����*��W_d�hӪ�F��8<�Ir�p[wf�:o`9�RI��$V��g����<){��i"~(ґ������Z_�����-�l��SH���7��Q&c륲Ȣ�Ai;q���W���{��oqp�T�]	��Ym)%�o�ӿ[�ZO��TB8�9o
C�\��zk^�7����y�@����٥R���/�F��u/��#��NA�N
eٲI�/Y�����d�
��B3�
��'�}7��p�~"Ih�1%.3`+���D� ��]٫���BXF�;�,;�,�����R�/�;��".�6"��ڊ���b�L���?�^66c��|��$o8�ҳ����^8"83�����,����i�o�q؇ڔ��}�|Φ���.�z:�ɽ_A�S��B�+T:�3��E�����8�M�[h�AJ A0�����}5�664��΂���xMZ+�X~���sQP�g�u[�X�=T��aE��_μ@v�I�g��Xi�F��� �#V�����^���ҷRDF7{�z���AF��˕�2-z��au\z��ӽ�6�����=�<�.�}d�fk��)�*�-��;�N��1�9�g��m3:����wHz�mE������!����O��yYu�B��˰�HV�ab'��J���6�T�5<?�Xv�_�(ZY�.x��<N�k��G&IPV?A��2eZ?�*�L��h��5
�V������"��͞3��p�� c.k�{x�l�H[�~���|�GPLY�P/
�H�/����b�!|!��Ps,'UF_I|G��q,�r�Q�.ʕG�UU�7�����`��u��^$U���BP�������K��9��p��1�:a� �j�=�@*e�;�R��˓��5i(���l]e��9B�cqC�$[�vy#7�U:��V�mM�n�D�"�h����#���ez�����	���7{����J�«����N��cG3Z��=���8�ș�����c���Vt��D���3�?�c�qج��-���MS�t�T��~Z��I&����$2L8K��p�7*6:3��:9~�k�X��3�꽹�$\�2�X�����ߐ=������57]��W�S���U��������6C�Aq|?�5�`t{��hF��=���v�dL�!���(��.�gg���J> �[A0ؔs�^�	j�vژ�pBz�[P�_/9-\l�ܲ�X���y�E0��0��.Ż�����~��y�����.�1������,p��8\�w��4Q$�f�U۹{��|��O�)�$�<L�&��q��̔�ԊM��'�!Cd� �w��H/��� -��b�H#�Hd5t$�zi�����Pχg~��w��=����y�vT�<{�35�eR�e~
m�;�Yp3��;m((���;9��~I�ϵiEyWW�%1Y�GU��1����@y+�H�@��CJ	�ȝ�F��3l_ө���EZ!��?����/��9��-�#��l%T�!fJ?v~^D��3��.���+:t�	魩�(�}���zU��p!)-ͯ��2	��] oALЍ��o�S3V�%'"�]�D���H��Y�>5iϝ���F��
�H𡸭�H�^�s�h���1��Z��_4�mN2���7x���@�E��E嬨�Z��� ��0stj���I�1�͖��?$c�|��j�l�	�;�I;%�P#z��gs>�n�D@�<A�h��G�C��q�ᇥ���ux���)*hԈ��춇G@�Nl�b�cԻ��_�a!t"Z)��������O��'rץXW��#]�{ߌ8 @ߠՄ�-�mr�Z<��X�YP��\�U��bBZ#-bFf)\���AQEųmGq�ⶒ*��H��Z;r����� �٣��:���r�b������6(�>��A>1�4Pb�`o�y��\kV�V�G�T�w#���Q��B#P�x.��q�Z�c���-Ex!�l�F��\w���⬩�8h�і�(u�J?���P��OO�F�c�)���r�̩���Ó�Lߥ�G?×L��S|�:��Յ��&�!o��hZ�V�r)����P��H�̙Or���{�
�
��8eq�U��b�?w�����y�vj�%�g���^���}O���]KKD�,�sW�� �ׂ/���z����kok�x��I���SD��iA�<	qmY���֋!��\Q��225t������O��m��"%���)���.rv����Ƅ-��#��ڹt�@9�~X����y�N{��O�Q˒*� ���[hd�Ŋ�|��~V]w~�A�}sϳ�!��ׂKP ��yfb%��\Î�ŝ렆V@[-,j�R����uŧ���C������4��YX [&�����	�=��z�@5l�c1���z�FC�n(�����i����[q>4�ޥ���ċ򿭷��uƺ�tїg�Qt.��\L#��%��U��'�}�G�����;�x��/��ݚ7����M����I�%��jG�&��5�֋���wBQp %"-�at���*���ɳ봭9��8R����y8��CcE'��85�]�����#��=��Wl�ŔY�^���I����`6?�o�lg1�����EEF��z��m�6�C�%�������_��RV�����*-�oo���>�l/z{�5�x�P�7�����o�ɴ~�������c6��＼�F������V�hi��-uh�&��Q�ه;����k���$6mK?�3�-T����� F�PJg���(Ǭ�ލ��yҘ����U?!e~"�cY�Tmv��g��06�����t;�&RN�6C�s�6�Kfj�I�Rs���#ىuh��6��P1
����K]{m��S���,��C�V�rNq#�<�Z����o�n����+����J�^���G����j����,���DObiC� �6�TU!~<2���zd�¥H~<��m�ڀv	�����^���Q,�dc{���|2cy'�������ש�~퐻<9����eqQ�67�i�=,�`5��И\T��V��������L���n�h������W���x9WսY�2���c�<�ϘlB���+�p?ft��6�#�D�����Ű���ҌZ$j�o�@,���ؚ[f��*~��d�a�f�H>b˨'�M}�.r����P7&0bl��l3�y�]����8B��4�1���p�6	�$�<����	���r�rs����~s�вhv�Fd>�������֧֭��}���Q�����6e�@t~`����L(����ؒ��5���bL�n�[{kQ���lf�n��ym�rp�֎f���\;99���(��l^ʞ���;�:��蟇�]J 𵻅^�AҚj��9T���8\�3�����'1Kj��J��	���&]�͂FQW����+�#ke���)��ogV&�B��th��c^!�����+��j� qww����N�����Awww���!����߿��p`�7����U�z�p�.�ۜ��x7%+B����T�K�������+)��(���^����n�b�w+n��=wmw��8}����bY^��!�YbI�o��3�������P� ��V{�Jj�v ל)pJa�nGQ��>��R�d<����,b(K�o����ܮ]	)��٥���.b�~w3��3]o���m��O��=f�WI+*�/���r>���$���"��N�d�"7�;vV�uŗ�z���a�V��=$��P�^B�?��Z�A��>P�Z7�+�Lϙ�8�;{����;�8�$�'`?���Q�_>�)��T�6k|���"S�kF���,<��Ltnĥ��4([C!}$�--�Vsxk��r�%�o;��ۃ��3Վ�i�n�1��&��'P�1�F��L��yfc���-N",.m^%v!�p�$f��F�}���kO7�(�+��YA�������k���S�e������]�Hiii������W..�PT0� ⮩�f�M8��� ���d���8x���)� %ā]�_�~�ӖQ�yv�[�BV��V���	M�-���o�x�D����lxPlu�����@JS��n�DPz�++H_���̙�M|}˫k2�}�D%����)�#�7I"�s'�;NF��)!�'K�IX=�/IB��م�Ӛ���QĂź���T���>p����.��K��( ��=���pmm-���Wc��C'D`l���G[�JT����Lh��7��/?�.|,�W�pF��`_ �D�>o�����0�4��M���#��7��zj�{�޵4%�)tdki�]�>�
���Er�d��:Ҥ�y��[Q[7T=�I��<^H�c���YC��8#�����,������"'�<Pj�B|V�~�Z��؛ӑM����F��x�8b;����P6��ï4v��H�V�y��Pa�---����u	!O��P����5-���I6X����-��yvV��e�!�QN9\�@��i�*Y�!|�QJ-����_���[�X�@T�T�`g�,^F�
,z���%FL�{}�=�W:��{s�l�d�r�a�n��تL<Ƽh�������#��b�����0H?��n]0y��eMt�i����7ڧљ���Ȥ�L~�3D��',�ۡ��n�k
��P���?<�W�6��iI����[Z���pp`�HΤ"�*+������P:[_)�& ����rx��%��￪����o�k��o�uF��PLMM�ă��h��tf+.��!���c�=N_^�ir&�����EH%��B>h�5��I0t�sA�=�u��DB�cB�qm.�/h�oũ�7��K���SsR}�^ę�U�c�Ѳ��А�u����uБ�����7u�V�������0Q bZ or- ����I2r9u5ҥ��sf���ë�����c	
���Y=�/^?4���F��]������F?5���j�U�����'��������tE��1!�K��J=t����M�eԯt��< �ZU�V�:��^$B�sև��L�[��@G�|E�|���/i��}�Η��_���*��JuA8x�T����(nN�/��y�S3\jX$Z ����e��i HD�V��Aa#��K�R���즥T���j�I��cj��sd�y?�&F���IJX_�'v�wU�W<�[rj�,KPLFl�i�a[{��j`H� �0�D+�X��n<�ʽ���"�d��k�O]y9��:���9�ȱ��n�v���T�r��_�x��_�����
�p��t�ܬ�d��<P�OQ�P5ăA5^yՈ�:�!ۇ���j��;p����{T���t���B߱�A��)�s�lo��r��Te�F ���b,h����r��Jħ����zT����:�� t��X��i#���&38�:ː�	�n�Eɐ=lp"�L�� �"��)4��=�����
c� ���A�6��[�1��m�����z�ֽ�{����.w�L���I��k���I5� M��T�������K|>I���d�	o�J���圁�c%C�Kio����y���N�����zF�W��Ӽ �!ˊ���8��<k0���<`����Q��ǖ5鉫R�D]����_!�s��[�8Ȝ/;������	<e���2��N�Jt�:a��V�&��+4��D������S�p�L!�έ�Ǽ�Z�G�Q�q�b^�0<.��2F������8na.�ta}nN9�,rwB���2�)J��5�g��Ks��كU/
Es;�q�k�4",�����%/9��ӗ�&�d�8�b��t��V��ݥ(_���{�K�B������j�,mP3�@��b��- 7KeFFщ��
Z�v�Ŝ��ضJ������!.�3�ʿ�iyԢb`g5� ������J��_�o�$E��L�׼"�[z�OUj�n����߫Ϙ�t"��I����%��;�Y�@u��KG�SOG�1ăVfNKF�SF��Կ�pȍ��Bf��Ahtn%Q��9���D
��R�:��X�]n������`$zm���|g����ؾ�q�K�̄��({��@�iY0F�$
��=�Zi3�qE�,L7���|7z���zј�f���c�znIL��3\F*�Z���9!#Z<n:n��9�9&〪9s��/I0�g.x�NȤx����*0e�b ޺�ĖT8�L��\A�ʈ�(�g0�������FA�Q�a	ѫ	�F���y�e����k<���ۨs����@]��㳻hA��$û��fdk���~���,����+S�R�4�:���M��ú"z02�q<�k�v�ʑ�H���U����p����iLI��Vj7�;���cI�bs7|5�?��*j�\j�ײ�T:�j��\͌L4̇�Q�N\������/��k�`;1�����4 �G�B�g"f����.@AVhͥs���r�=���G�?ت2����S�x"$���h<$��Os|��nQ�{ �x��Kg5�b��D�ڬД��xJׇ�1"M�C�ʬ_��]c�T���`�V\ōy����*B���9+�dqW��KR<�i������r]x4Uw��k��}�FNb��%�qt:6|*��P�{�O�s|�LP,�� FƉQ�La�y�&U-��u���@���Ȅ���p�n^]G��&{VZ02J�%�)(0Qc�:fb�ķ���@�i7V���3�u��q1��\zؾn�Q{\�T��b�Ϣ?P��8�܈#�D����˿�W�����u�tu�S�B�i%D�l����P~�Kt	�iRF� D�1�-):0|� dpa�a��w�U]W,l!�<���
��F�H2��U.��,�r7u���.I�c���,�pV�"G�ee0)0��GA��Da�|����Ad�%����r�dɄ3��p#�#㇀&��
o��1��[^���U
�f���c0�)�L�A�ą�de�(�ŉ5�~�CG�Gxf�Z�#��r�D���ķ�F�S�N��jG>f$S�WF�TP����a�_W4I�*�׻j:�yA������`�j� t�$F�1�Z��ʣ��x�����8M���g�M)e�e�sHR�Jit��cR�� h@����Kz�u%��+���� !�����b >��H��(�`-\D�b0*�(yT��1&������a�����.c��7���v,_4�"�����߽�ĉ0)'d�h��_������H����R���~��=�+��H��T�	��4�~DZ���3�F�����뿘��z��H����{%0�1Za�p�t_OЇr�>g"�[�6�K.�*���+�FNl����q���k(5��F.�豮%�0'��f��Β���&�C����G��p9g�`5̨�gnFR�	��(���;U&}>G����1h�	����tp�b��!2��3�v�x���G��ߡN?�P�-|�ߙhK@;� ��33��<6V<Q�#�_Q	�8QX2�e��%ѝ/V� X>�:�+����o�6h�Nk�=F�YnFt�AKC�i�J����ލ&��Z����rRG�x0��*Ng�ܛk����� <M��P~M@��+�\q0j]�jG\A��=HDv9l����-�m��i;ziZ&GT)�;n.*g۝�ߓ4�ɐ�(���D���	��D��|�E�o�"���C�՜"��)��NF��|�q�|3Q{�(��=�q,X��\�f�s#S���}�MW�	]�:�zO��ޜ�Z�����A4$j�%u��wPh���U�������J?�'�*XPvH�Z�H�̱Mw���L�V�� �&��F��K�*Z�x�j*T�o_ݥ?������cO��
?(т�^6ph���5B�W8"~ȬI�'P�<o��ʱ~3M��)���؃ �1۠|5M #�n�r1��k0B�W(�x]�χJ�Z�͟��p�v0t������� �}��H�Zi�����=H��=>�( �tQ�lCX�W^�����L�d�gb]R%��i���}��O�d��Wa
;����Z&���1/^)��kBD$�N����Iq��gߐ�ˢ:�{�=M����&���%%�����4���9޶M�(8YZ�Zb;�|1�9hfv�G,}���4�<i�ѐ����m~]��M�g�oĕ!^}^e�%Q��$��z�!Ѽ�&G��,��H���F�
K��ϻ�)s��HO_H�3~��c��bj��̛`�]��	Vz|
B�����t%b��詫Q�������ҏZ�b����g6ܒ@�i�=�I<$u��X	��v�R�6��Y��
S����%�O�Jԋ�
��g�/��|��]�/�g\m�I�Rc؟�YJԋ�@��!�؍;�E~���i��L!ar����,��x�o�7�E8r���<6">]��_�BS��&�	6�w����Q��]e�E���Ѩ�E��������� �H��������m1<����ƺ[���Ӥe�g��	�� Z�d���$2
�J���Ot ��NCTj%��,g {P�ɤ�Xs���Y��A��\����Ru �`����˕��/cGI�tE�f�TE��A8:��*Q6�y+�|����P�j�q@�\n7���P�J.v"�k����v�R�p�D�Q&���hMoQ.��fQ9�X�M)rتt$S"�n2��$��եwmSm�Q-)�^G㾌nl��4X l6�ئ�l]=�����rbS*�S���)�#���8���-�x�qkS��~vFj��t��(�fl�v�6�y,�b:���f00�X�,�k�XLţş@<6 KE�&��6E��hOe��z݅�	��̟���<MF���T�V�y��)�%�5$�����u��Q�k�D�	o&�����.=�p ��@��PIϞ
E�i�P�U?�&��2��S�U ��!����<�� O�q �Te�wlᖽ�ܙ�״���>0�u��g=��ns��BP��D�OB��|����<��*�@'��݉f"�A��t���+\�6��뤦LCm]M!ߐ(�35���2,�MT�������VL��?3������S�YI �G�_>�f�76� j�K�� �3�DW�L+a���C�q��,=$����_߻Q�Veqb"��k������n@o<��7e�$f���~�'��I�tN�	$��D���޾没��}r`��&�1tR($q����-*�����0(�G㏃�d�Q?$\���7X5Y���؇��fm!L�8	~�\��9V��Da~f�� L����ig�s����=���x� �84x8R��.�*�O'�OP��_M��HK���^u��x���x���L��X��1ߥϚ��$ܻ��wާ�ʧU�[]�T̎��j�G�u�z
�E��3v���9igeW����5����z=��������n$�X��N��8d�kqOqH�����m%�|,{F�������'�c���[�)n�]�Wm�Z·� FN!-_���X2�|pdCu�ob^��}�RfDy�>j� �JX5�\����*Q�Z��?��"�|��^ �:w�~�~�z�s�|D'Gf<剜i�����z�6�y[����6�"tw��p*�D8����y;E{��~'��ZC��̮Y׍�=C��U��ˢe'닮��ʯ����"��A���$� ��{~D��	Xr�8�L�\`�S�̎�c�؊�Gg��<̊����P� flL�jʹ���*��Oµa��+OȈ��T>=�±S���Ny�:��[��X����~�yC7><��{�h���:�2��26웈�Yk�x�W���l��j���N#v���=bܾ_1��wR���۟�S\k���||L��o��I���v�/���j�{ ����z>�,���D ���e'�v�G\8`k+�(�P��'��h0�W�+̤�j�*�qêSu�h�cu13*�D:�N'Z��!���A��E`���O�5C%���Ꟙ�{�z���Y&���P����?���wF=�o[n��7Y�p5ԓ�U���`��b�_F�U[�`��3ǩ<M��f8��](��c2r@t �0����.N��X_��_�Î�*����Nn��ȇX�ݜ��Y�������&�P�S��u;���s�I�k ,8ks)j���������}� i�~#o�g��~�4��]{=�*�Ki� �!8����=�1b��}�1Sg�2U+P2��L�˿C�5��`vu��� Zv8"T[�r%qW˝�D5L���D'�4�~6�,<T%�\D^^�h��o�1��#)w&�*jl#}%�����rp�XA������O^>�����y��ŤL�e�B���#}����2�=�}<��eḦp����A�Їf?\թC��0���4��3�-zN�o�Xy���rw��e��D�нM�#w����{m���_%�I��%���j5�}��)�9���6abT���vD'�i%A��0��k%}�wT��Ɗ͉���W� ���)dF������4�t��� W�0�=�Jj�\�,-G�Կ�Z	~�2�Q���P�P�iX$̧5�E$�8�b�R��1�7eh\r�+�!g���}�8�429x\˦�x[~�E��I�ؾ�g��8��`�������ha^7bFvqI��;:�0���N�lޱ^�o��?Еh(R��L��ȫ35C�t{�����I��+I�0zu9qII�²�-�e��fh1��H��`֩�d,�����_m��((ŵ�|p��ߙǧ��� ����Vx���[�����	[��b�������+W��ܨba)��A[�^�۸8�Z�"�������Xm��*B}�3Rb���y��z!N�B����%�)ma$��Cp���8g�\��(����'Vk���R	��k��R�y|��#(�$j4�Z�_�N�9)}}�;�+�#;��y(�Z�7`�%~�m�4y�Q�ɳ:K��\(��ݳ��!�H�6�}�ǚ��X`����.�G��1����׻ƒM��	��0!5?Tt$/7�eև2ɋ+jTd&&�y�ާ���5�gw�h{`�݅�\m�l@�T�:����Z�U�HIea���3;�M"����tеƏՌkQ��L�0*��1�6�"+q5H,�	f��ě��:7h��iE��η4;'���\���C`m<���T��%35gx�h�B<�d�P�i�lm�\�y�� KI��Et咿P�"A���l�2�t�����im9�J�`��6�߈y'_ڹS0@�-���7QRhԻP�\^د^�v�f"�>�a$u��-�	�[�[9G=���Z�=a��Ɏ���L�2���C�ZX�G�`�	���@�1���Y�K���S���������t�.���2�8FM��N��g�#�5^.��ِH���S0�*�ϯD��N�H2��ޯ&y����q��z�]%���򢍮�M<�Se����YJ
�;���
���V���g�k�1���_w9o#����߶"�>�/Mt��$�	q��F�|`�W<Y���s�34\��7���6��]���W�Xъ������HH�^�*5��C�ܭ�2���	iB~7m��N�Y�$��E��j��so�P"j܇�K�Z��ԩ���̣�`3gy�ܶK��� �� �ъ�6��g+0���o���t���'> 7�c��Su�����:��CƯ�������_�}V_���Hv�Db�䇪�lu9+�lXN>ZyE"Q�|�$6P��HBl� .���bwN�Xj�'	}���Fo>�]�:�/1qM�Bc�1=AX����l�~��
��N��wu��e�b�ԏ"e�}��n�,�5�� n��b���nwt*�(2���e��/ԅ�
�f��)�i�;�{�60�·��[+��?<6F?���o�~�ɫw2���޵�A�)KA���e��S��_R.#p��6���` �'?Iۦ}�.3�'�;!�"i��_��;�/fq����9E'ey�d�Fr��!�e�S_�D��@�����zW�ER�{>�).)u���u�B�*��w�������[?�����6;ﾛ	�o�����&s��>I��(�M��B��A��~M<D�↦�bq�W$�N�������<�j��M?��,�m����|\��G�OV'ey�[v&�p!$�r8��5�0g�����䣫�����L�P��cl��nv�;���}B��p'h5��C���ˊ@���R�j��O�|4���Z��xL��xx����^�t���.�`3Z��IȦ�.rsRI(
σQ���ri��;����1KfH5�uFEB2�̠w#:4xg����Y|��fJ'�j����&�h�����e�.T���D�.2�x���a�u�%q������fH���D�G��\�'�#�� ���+�+׻���_v-B�Eļ����k�[]v_���9���-��m�*Óf�׳�%��K��Z��ݰoy&�N S�n2g���<R�/4�]['��v:�q#`�?��L�*؎<	����V?hs�4%z{��t���}����eQ����)�;O�>�zbR[O+Ҫi��3=�9z�u?J��d-�AR�W+�,<ؖ����9Ӱ'���Q�Y��9�b��?Y���
��	�'��Đy��Y�v}�X��',b��o�x��p]��	�O��X�ҟQZ-y����<ʵycxU�T(@A�0h)�����0�@yh-[����%D3�V�r���3HP���S��ŷE��#��FtϾ�;!L*,��m&U�i;� +�B<� /��H?�l�`�Y�K����p��8�=���v�Z
�b��mt�&��O��Y���r���]?�1��o�w���l��ؐp����L��V`��d��%餓�&�������T?.$�z�F0C��e�by��p��$���F_�X%ϙ�����������	�?5���ml�z�������xU��~�������ȼ��u����g�����ޥ
�,f����jsU"o}�LGٓ}�^�X�P�x���hM�0�4B �cS1��o�s���ݐ��sd%��Yzl�ģ���9�*`�kj�kNU9<]	�u}��o��B=�+>z�Fr��_l0�v� ,�y]�?�Ѷ�wm��-!쌡Y��[����3��������B���t3�K7���#�� !-ºK!�#8�s�*���Jp�ۗ��dO�a[��[���" ������ǄşC�yQ
��<#������X�����I9-�ܘ+��Ȇ.Wz������D��H�N�7HZDW-QK0�.̊O>ϻ���Pt�Ȑ��B\6z�՘�D|po	�X�'J)Ϭ��1�svTӣV腀~��K���S�NB�83q�zJ�ז��گ�á��r�o�Q���hͧ�|&��0@��S�j���|�{�\'���Y� _9�B�O�P����+���[Ԟ��gš�u��BT}_� �J��A���O�X/��)�p
X��% ݂�	�� �B��
ε�8�s�gF�I"�S�j�w��j�q��?�E�(7kOO�1�m��`m-���K��<=�ѣ�t,��8��?n�zQ�Zʙq�ˌx��A��z���=�E�H� r�[�(t�7��V��K�M_��P��(��ة ��c���x����$L!�D�j/������#��'!킣]�]R0��^9H�*l���ӽ(�F%��'�:��֭�Rf�C�r���4@F�S�_>>��BtU��t�s�Dwe�ި%�������T�!	�d�3sm	���(z�?�G���R����z?X>��0E����6��7����C[�;0��u�����=����Pb2�����1e;> x���p՝��Ƚ1f�q%��p����'ȫ��b'�J��	�>F$/�Fm���P�ˑq�_����HQ�A�i��V.�]�-?�*�r���Q5�����a���c�K v��^��~DS#;�/��(��~�����Ϝ���&e������\��R���݋����^�z����jOvS�F�]h��-a*/��T�J�eFc
N���~/ˑ~�Z%�s1�L��/(R�í���н��Q\���ҝ�u�uT��ܷ P�;1�=|��5�U�L2b��{L��$������!.9���!+(���Z�R�� N�-��S�`�[���^N�;L,8S�\X��s��0�JG#(t��ޜ��ޗ0C��O��$<���\]5u!��i��=)%��L�͹�:��z�t6w(lW�b�Yn{52�L�f�4����
�.�8�ղ;��g �:f�d���r�m�o�V�ݜ�'�	����:���6_�\i
�����b]p�~
 ���;j��,.�������f�S��b�\u��:����Nl}��[��tE��jČ�{/�f8��)b��EA&���@ļT6�axXퟔ6� aRvgjtV�H&�+�K3o;!��Nkz�1����Tk����oN�P����7���uIl�,����̮�i8{z��K�'�U��y�/����,|E7z������zp"�?��z�U���k���|֞wBp�23y��� ɶF�2�(x�N�[�@B��LM�-�K����4!2�����e�h�W����G{پ2�ha\kĎ_T�Mힻ���d�X�7t$�́�__�c�rÚ��P����ƀ7��Yϓ��y�0|�> ��a -�s_��ȭ��b]݂S葩��|81B��C�5����֤:>�K��,GR;>�6/d'�E���(�|�T���^7���{:+����L}�i�.���ʟ̸VF����{�"��v	��_]�z�~K��Z�){ի+Q��'A||���l�/�2�D�9��'H�;��;���`4q������p.���$:V�ʫ.�� ԝ=�pei����i3�m�L���JHAǞ��K~�ֻ� �����,��T4OD�N"ʹ*V���5q��/z2�+�����TO��D����}F
6�I���/������l��p�D�4W�Xѳw�{V0t�|�E3 ��ٺ��]�D�<��g7�I�(V2|�z�[���m���M� FӼ�д\�]�}%5�N��ams����֓��?����r�E���k�#x^�<�5����
ѧ�4�"8��^u�l�����4]H�$.��Y�?�ŌUNT�r�IEq����Y���}�n k�<�����^�W	�w��ED"x��-��ʬ�����K���ZV1oj�0=;�{�����Qz�͚R�c%�ps��VX��5��L�W��L�i��������D�rP�R�3��&��]&|������b�HQML�0#Em�p�zԩ)���Д&m�Ek��B�)V$Sv|7��iҸ԰]i٨�aI���p�D�&0J;��>�P�ɂ?wo`�-��?��|���?O>��R�y���>#���L|�Q�D+���ei���.^$t{��&.S�֛b�;A��`��#YƷc���A\�8���7njp`O��ֻ���9�H�]�O-*ϯ�a�Ajj�#b��������@i�۰R�`�Ǫ�i��˭Xy��
��@D禉c�1C�ޘ�m�+��[� �ǫ���CTw�x?���i�AK�~*��02�3����T�Ԍf͡}��tz]&��ސ �h�n�}�J=8�;-mF& Rc���B�H@<�1�,uGS�O�c�E� �6��Ƌ�tN4��{�.Q``��z�iP�Tfjڮg��JKd�ع���u^.�t;�y2����4��e�A�u\/������3a3a@�I�b��V��Q�2�=�{���������f�>����`��[~s%�[�,�//0���V��~X�8X�v"|�a�*ணf��_��6�	Z�HZdqrO�?�n�-�I�w��6�/u��!�6�j��е�	�J{ �q=-�L�B��t�W��;n#��f�y�rÿ���ĿR�T��v�ۮm��O��=)�R�PN^�������f����z-��nC���B^��0���#����Ķ	e������שW�j�e�uX$�[�s�ß�S'��g� ����<��02e߇_��/��YA�HA���b�
� ��O+=����LȞ��-52`�T,n٭f�_tb$��!���}~�����l�LQ���9y��݆fDp� �]:?��}M���Ǒ`1�^[5���\P�bu��Aч��A,�s��7�#N�7G���52|7��<=}S��i4(�D�K]F�\����9�=���YyT�<~)��ft�>�ּ�,0J��y�Zp���@��.��ΉgS��R���:&��C��+���`���"d��*��d`C�'�]\��}`P`���� ��*NA��hj����E܊���ٓ���@
�nm��J��%s�Au&�%WD��3��Z������BB�{��V|H���i[8z�k�	#���w}��]ZW�b��G:�Bݭ�R%��������JB2֑P��~E���P9������\�d�������E�b��)���g;Wq2���6�=$-5��w+^O��R�%�Oi�^��$ϕF�y����:D?Vi@h�bi��o�P"���t��� �n��=9�{�d6fZ������i�o}cԦZ��~@��\��v�����#�%,��x��Ɵ�����9S�O����`�aV�O�tBw���y��Ƞ(q��"����"O"�?�[�p�p�RF��gC3`f��#��F,O�K%4pp�>��y1�)8��
����+��o���غ���8Ko�8V����}�r �J��L��,>3W��Fd�K�E��Mf�Q�R���١��nt���E�"p:(�-9�Rb�M��h,qU�$F����_����%��"��[ӽ�����4k�ղ��%g4Ӓ�tp�Dj�rs��	�aT��T��'4m1����`�+�48c<?���2��`f4#B��kJwhnw�X�[M�!�fsԃv9�k	�ԂA���EV���[=�:���Aiɨ�TdA�N*b!�~
�:�Zu�H�b@���=dZ�EJJ��YDƀ������ᚷ�s��!�g���[w,�f�D*����qU*E7�cAi�����4�=���������Ax��uw�4 &�^�'�Q��]Niu�ƈd\��NS��ɀfo��*��?Z�T��]�r8�OlW�f��̬�_�ޜ7�fP�c��ҧ|^5�?Z��(ˇe`	Nu}�cp�`A�V���7v�ӑ��yi.r��b�\9n'�AV�j�-�\1�n\���J�"�
e��?�����ÿ��#S�)��kdWb"�c�i1��d܄E����.r06��feܯR��V�ǯ�k�����W֥��L�î�[j`����#˘��HJ�����������=!�'��w��5ր� d��׹����U-�&M��\��=P\_�9zijf�-�{��U���(�Ug�mX�v�s�)���q!u��	�l�p�߳uW�8��� J9��ND{I�=���BhJh%�j�m2{�~\�5(rzӎ���PfG�њ/�W{��/@��0$��q�!��n�͞5���CyƏI�������na֤��P��_N`C����=�U01Ћھٮ���ô
��f$�:��P�k��I��Vg��7���E�dQ0����[)�y�z9�A�v�$�j�w���Ǉ�&r�+#����V�G?����'�B)���OQq:�LBr�E}������`K`��1��z<��HPe#����Պ���Qr��g���8x�x�[�Y�4�d�E�`��.���L�c�����ّQ�d7�jN�CL�	)����e������kM#�^@���J,��K���o0�e����wEy ����}�q�������iI�|��h�������2�(�����6O{-@T3q����7��۷yu#~��j�,`4�Y;�m	�cϷ�v�Bm��8���%��%�A���qo������B�@P����vs�B���h.��@�ˎ3�=`)Ӄ�;x�lk��QɅ�OK��I�/����n^L�����ӵ(�ʝ�b�V�*(6n�q��bb"�W08�ޙ�>n�zj��N62����f0_��A���UE���r��W?��y��v��{&}�`b�Y���b.���,����9p�(� q��~�jdl����o�b��BX�1�OE����Y��v���?��Kٷ��P�b��&(&U=��)u_�_��6h�]���4ႀܾ�U�:$�G{���GYNK�q�j��CP�����X��!�k�_�p��"&�N�*����9�n�#�G nq@=��J+x^�$�<8����SD�x�ޝ��@E���0��e͞�v�ev�<�i��ܫ��|��kb��T���xn���^9�Z�����7󀨟D���d�w�Z���\H�US�4곁�!JbC��[z��^7o�;�{�旞O����}��|�<���3Ç��a�P��fo��a1���c��6ҹ޿#�C�,Ȫp���A���h��.��J'G��)B�S
<\nj�¹��k%j�.s��4��5�}�,Ȝ�B���t�F��"?�0�vW?Nf_I�?��m	:�7aU�z)����thI���\7�޾�T��׋��
?��V7�$�z����ɭ�觊�����
}�S������4P�H��+�o^-w��D�!�Q��V��Pߺ�>@�⺖����s�ϰ�e�g�%��'����=�j�ζg��fďsˉzW Y*��1�>$f Dx��{�q᎘�
s�FKk��a�B�F�aO	�G���n���F��>���0gEx\�;�����]���i�[6ˠK�4��8���;H"���~���MP�%OH����M�Cf��o� ��s6��yq&�j�T歫[��^��A�3�KSS�^׆�HgӨ�4ԃl<���y�Gfmχ�=H���&� ��2j���A�X���z+(��͇<�èb�)x=bth��$R]��# io����m*3I����0�NPz�>=��4D{��3���(g��`���!�Q'G��5�W�_��|��	%Q�#���5�n��D��R㮪�t��-E�W��?�M7�C3> �Bn�
Oy�U\�9�ָ�L�Ń�jm�b��)D��.LT���Ί�=G�A!��'f�#�O^��Ԥ������7zҸ����+Ϻ���r��-�Y�"zk�z}>�5�a��3����뤔F/B8*��!�2�H��u�@�iOd6��Տ��߾�MN9
�+?�etJ��4���;��w�/�J$b|�׏:m�C���MyX+_�鮳�-�B��7w��	�J`��\���uw�Q��(�-߷�ک�+n���G�]Q�� �����
�9Tɑ���YY�^kKѸ!��i������6�'R~�
�Vb~��:��fAD �<z|(�z����T�	-���๦��Q��}L�of���T��fmgm��b���3�G�`8.,�=��ż���쳿� ��rŤS]��D&}>�϶�ܗk�R�k���Ee�{�,���Wv����[�6��U��:��wu.ln̯��-�>f�8���^�ػ9z��pJ��Sz��ݍ� ��	<�.����'�Q�����j�E�J�v&ɥmw�A�ef(0FB!�ڜ������u�m��mz��Dڴ)�3�������~s6(��b�*Zp�,�v�3� 6�``���$`���Da�d�2>z��?K�������dI�e�\!&�vʵ~<���3\Àh��t����)���oO��*⎬nO��z}���$��=�]�z8�OU��)�Nأus�!��
:	�=8���u����)����\��`��<��1��r��4R��Z�{����W ��4�^ �������!������	��w�<��v�|�{�
�����鞖sfzz�	�|w�mw�.��wZ=6�� �ջ��h�<r�x�D<n�͸��^�����\����=C&�vs�rȲ�#�[��߫�X�����u�.X�a}<�h(�/�	+%�q��F�֖1�U����	ފ��!T�\I����.`'D�ڶV�s�3��y��i!*���DL�B�#շy��������1d�M/�$�4�8l�{��&O�f�RR��{�z��wf����'�n��k�����������{j�9їӎZI}�S�˳[M������q5E5K�:�A
��sdwǪ_ie%+�W��0�5�"F*믖��և�H���s����_��-�8ǜ�~��`c+@��7��x������B���Z�8�m���j	�wv�q�!�� ���æY����|�1@dc���$�G��t�B�{PCSPɏw���4�BJ��C��җw��r�Ը>�5F�㺫V^>�G�6lY�l��@M�?D��kえ���>:�/I���Y����pp�K&�����w���0̍[We밚��:𮦗���.Α�\�v�� �TZnY �#�]�&eL����H�A���x�x�y��N[��h'�E��V�Zb���-D����|���x��	���\I:Ǚ3��SC��h]u�%�^3�n�u����#A�Y-G¯�s�����Z݁�����5�ߔ C7���$�~�C��!`�42�o<�!�Dvmr�dXP���y+���:��O��RT�Џ��hh5��x�VeKh!߶�o8Hi�Aꕘ�n��.�qfK��K��^��d]�Jt���`;��AO_9�e7M�4�s�Q@&�׽�L���7^��1J����:����%8^ RS��������{a/������W~����#��6���&M���mY۽|ޓF��I��E8���^�e�e���#x����ߴ]}ᐩ��
��#ף�������N�x���0��C�o���!A�M
�m ���]����>u�?:��zD��q�� ��֯]$
�������������ý/�P#�0֜�l���yno��q�8�GE�E1bE���K�D�5u^؈����9I.����P�D�����A�}:�Q�<~��8��l���k����k��J�if6*�Y3���>H�JZL�#kc�������R�F8�0��$]]]u˧@��i~��=w��x2�̃{�K��wM�9�^m�����.��]�y�/犞"}�̍�v4)�"
��.S5�˔O-�&ժ0ҥ5%o4	��9V�CYhw��KC>�Ee�gc΢5N[}���=q,Z�z`"��h:�
�J�ݽ�ܽ&8���:�`#~>ݎ>RQ^�C�A�ʿ��ڬ���5�o�E���fg^caipL�:�7'�Vwvv
h���n9�ӕ������<�~y��4>az
0S�pRo���(�/)�b����m��I�0�L����5T+H��z�>VĚ�$-��kXdו��!rm�T9bZ�������? �{S����+�l}� �tP��Aj�d$�sa̕�&5Q�3�&鶵��3b��|�죘�jS]�7���9eH�,t_��ٷ�J͛[r�QD�����C�lXp(�w񉉉����;��zY���!?��OQn�A%�
��YY��3���dd'�F�괫eddP}	��f�����Dx�C�l_�޴[��b_�2�@�3+A���YCz�?�X�.k�G�?&Y��`D�؟�L���+nٱ*J]�����q��١B6s�/MT�Q]�I��*D��"|e)��%�#�r�WQ;rC-,[؊j��a�<7wwwS�Y�OxH�E��E�$]D�?�c�>L��V��oʗsF��L���zvnH�W�"r���@���<lדwu��/:�����J�ێ	�q����*�^ ��;�+8��/k�̓�j��Rr�]V�$z?��qD�uB)�<?�d� �^SZ��A	'Dnjl݃�ˋJln+"Ȑ+�4c�P6[*#�kf[�q��j��9ǽ�#�$�N��0�*��vP��x�6AH� 9K�	�ώd��xˀ�'�O��,�Hn�~�p:�9dn)7����5��_�2>i����\�d������<����o�7��9@�y���f�T�<VS�8�By�rP��d��ረ�o�UPQ3��B�a�0���͔+�p�ڎ<��+i��zA�YdA-�-ftH���&�*O���T�˖�7�d��O��GJ]��5wx�ЮI�.}�B��Wuy�^81o7|LT��D��ϼ�l�^'ދK�d�`��X�� ��)cy�,��"f��IL�֥�xgAo+�2Ej����[}K�3����T,���W��T���c届�vc(�	���(�햙MS�K9�廻@���~.2c)�����=K>t�>`�q'�d��O���.C��H*OeZ9�>Am�}�y�{X�"Չ�������uC�廂wN*m�JN8@~��X��bE�$�����a�%�
%[t�0 �(@�ӫ�5�U@7�
T�|z_��/��rY�1	1�kq���}�7����������R������ɘ�t3#���٢���ྍ��MT��:�^�a�:�2��"�ܞWu�7��/�3/;h��a��|9�טL��k�$��ׄ�j�R��G��c�~
v��L�Y�t�p�Ƹ�E�۷<} 9��{-���]�L�A���N�d��++�`g�h���X��#�t쵼��du�.P�� �xb�`�S��H�%;�&H�<,��Tds~G�#D�bF��v��ho�R��}�@m''��'��?<� �#�+X%Xg��r�(?;���ճr���jw�V�²O�q�w�MTE˂?UG�(�"h�.��[�����;�N0!}�J�G�,1/��^AbІ���˿�8���a��e�FY�3���;���܃���J��s\�����v|{����n�(-�1x/��V7�l���
��?��@��}��7�����M]Zk�[I{���x/��KvT_s�	���O�1>S��9�*=Ls��>Ϟ��[�EO���_(�v���#�2q�/��}Eh���Po�N��ozJ�+�(|~?%���'�c���~�g�V�o�9�:���#w���O����-�"��sB�5M�j����G�b��w�`"L����[ȶ]5���.Zs�'F���ԅA"5�zUhuϧ��;ᬿեA�9`�ć	-�Ԇ�l��1���.�5�Րy����삭��������L�B )N�7���Wo.e��^���)'=�h�D�k4��s»�c.h-�����ףc���h�H�l�#
��
�~=���1ӈ�_��-N.�zD�7��It����t�cQ�
 �$!eE���:��B��bcʈ�nM�(n �$
��uZ���l^;`�2�{�wez;`>�����]�F~+��_�*E�r^�xF/���\;lx�N�G7�7���I�ȸ���%�U����C��pe��KC��G��3��?
L6�#=�ʶ!������:bh�?��F�	0?gZ>{ĵ�ckK�g�c]",�l~ $��Y�wl�ԾX<�vh߮��5���dh��0A���MS�L\I���׵?R ��&-9@���3�Ƕ5aXvN3՚P?���~/�2/�]���̟�މ��.ӴQ?�v/���H��/GyԌ�r>��VjZ�%��}&����y���X�-|�x���I~��,��mЕI���g6xHxq�a�<Ȋe��n+������1^[�떵���b[k��a #d�����3ɪ�d��X�+灟�,��]�GO�j���\��/8O:���Ž��l��$�r�_)�:����A��>����>oTOM3�Ŷճ`�Xc^m�Uk0=۽9=[)I���w2��a\�O�C?�Cn##��_��c �U�V��Ύ��E�ыv^͏�F��0hq�}��
q�:>��:��,��L��(�^u�[�P�(B`�GW�"��D�7�v�f8�#$F����h��߶	�
jT+
�i����<;V�t�r��ʵ&��y��+��R�|�3����m�3��k6���L�%�C��������T����3&�}��A �7�N�;�8�hԓ�i�P=K��S���?�4����Lc���'D�V���N=���~��4e[�xV�J	2�܄�`�n� ���e�k�?�?sj��.].^k��tğ�v `A�?N=I*��k"��(�1k�SE��R�B�d��9�\d����@�8	�-��q4��	'<m_|c���Z��|�}�}3\�X������ D�i@��a�W'ǚ�od�����A��ALB31+�Is�(�uׂ���CX����� q�GD�bע!j��G�z�J�|gΞ#�T,���'���u6)�EQ!��VB�Y�ߋĪg�O�KQ:!�X15���(oY��FՓ h>�9���]zy�sSɴ�Y�37� `z	�X�)EX͛^ZLN�\Wt�lV��6�}�/:��c���I�w�����:2nL�èȸi��ʷ6A��%����i��e���Y��_���[�u,�'�M�Qr���V�)Wh0�nk�6���&�׋#ߘX�H��жY|��`hB*��j�RFp����d�Y�Ż�"���'����Hg,�7�-��N%yn�S "ol���{o�F�8b]���j=�N��Մ(���[!��|?p�F����Cl�b��@��NBX��B��=M�.A$@�'Y��ķ#O�(�8F��le��`k@�G�V�:?BR|��.�5>����Ӯ�`�;˲c�&?留8|���n�=�k;�Y�=���`Iаk}ۊ����9x)q���_���$��rP�TU�H�/��RO���~đ�z8	� aӁue�ܡA_�r&�g�J��ܣ����"1
LU<�Sۉ�5��˶��,j� ��8�<��{S����Z��Sκ,(!P��兮��b
�FV���Q#� �
,�W�8������v���(����_�������x����p���Z����"��[e�?,��}����_�9�FM� �2�>�T @�1��a�Ι�=�π���(��@��8��	#��A��P�p�|(�����sA��|��S�� .2��OV�s����P���
�>�P1W]����?Γ���l���U����cX�U�C���J%6L��3���a�f}W���;�&�`:��]�eYX��ri%i��>;m�8��vM�T�����2<�����<�暿���3c����M��H�<��@�&�}�\�ĭI8N�����D>�A��S��PA���I\���6m
s�gO;���z�h?>�KCJ^���\w�L=���\����Q�{��؟f�t�;� ��(���\��~k} �kM��ٸsQЖ������p7�*��9J�y��[������
P���Qf��Q>��ki��R��1�h�d���"Ku4�[�5����G ���Mc��ŋ1^�x�&7��,�DwNFF�y+_Hf�%Ƣ��[��q�j�����V-�Y��;�1'ry�?6�x�����&�Wҩ�"#�Ĝ���
�T�U�Ek��ï�'�������ul�_G������D�0ṕkD7]����_������3�Y#x���Ċ��d_������*���!�X�_���aZ<�8�Y����9&V�9�Kz����VW�O���z�kj��ϿԂ���m$�޺?D,����f�{�uۜh�P�}ݼ�╨N��>�RWjK�n^i�w�YW�H�'�	�\��i��"4���`����N&�e*A��B� 2'%�L���:��_�����s����1)�+�_~�nl5��|D�7�^�E��p�4]W�`EGm���eԑ�{�f��Wt�f?!{��>ߗPi��h��q��fX��v��v��j��e�)�w@��S�O~p��m�b$�+�i�>��%. �@�2Ղ�=���A���v�vK�"��&��Z���$�2�:ؘ�*ĬK-��Q��[7�#N���>���Q.4��q��]��ޢ�!�����Kf�l��p�o��0�,�� �E��v��/��}%�Vޏ�ȃ[Q��_��PUb?�s�g�\���e��.$�?BX�1?�m�|]"�3!�R0�TR��K�iBC�eHX_f_j!�!�J�l`��8���L����Gs���qc�oxQ֬�N��\�y���Nx�j�`��r+p�fj�t��H��$�zPGA�T�8��;���Z�B���}㤬3	K�n�#�ݮ�X�l�MC&��������H	�����}�+q/�Hx���-q���Ce<+�X��2�����n�&Ѣ6G��2�5�ח7k�9��C�ͩ����ɐ��/����*��Yh�۽�o4Kh�"1B���7�LGp?���z?o6���ح�И���q���F�dxm���`3��q�Z�R�:����"����~{Du�[#�P�#2?{�_�*��AnѶMxS�H"�Z�B��C�&�?��S�b5�D���>���WQW�[uLXiC�������<Ն-O	$��/F�՟P|�kA��e
Ҹ�M��]����x橆b�T��C���021:���-�����Ao2jc�
�`bR~`X��+N�N���H|*�@�o�ݜw�:2:�vlV��d��l�k�@=!f�G26I�QX�/Jra�����{6�4QF���^�����G>W"G0zs�qn|�t�C"�/"�1ˁ�`6y��6�����.,��[#�Z��D�����>��5UQ�ذ��-e���l[+S^�|���A\bLπ�P����S�O�5��Rrz�_6's?���jAp~�é���cC��7Y�mCU
�Gd|٬�/~O��ي�D��aˋ����CH����J=������W5�E�f8����n�ѱ������)���ֲ�w��*�A��'qQ�w�����R�x�h��#?�~�7n�����ٺn
4=&(�̓T��O�!NnRh�ciƀ��X��ÃKP�h��Ԃ�Ǆ��"�<A-�DФ���g1���%b�1D��i�����b�[���)~ݸ��	 ��o���R%��اv��?��s�����]dJ���g0�y�/�>�R�&'���c]�+���fx��j�����2�pq��q��%贪}Ra��H�ӿ���S/��[#j1'N���`Ǿ�:<L{8

�>$�����fzW�p�:x����8��\"�Xbo�%E�/�qz)�-[�Gp����6����FeR�ì����Z����'�YK\1��n
�����͜"|���p�p�=˫��~�Xz}Q&�	�m�dx��hL}zq��3{��빞:fPy��h�U��y�ӛ�i��W�!�b<�.{J�Uٜo'��(ة@��)�(�i�i)Χ�z)�zb�3�5��D=1����n��>�/��j�����f����M"Rg����	��Fi���d� � ��L�����SM%�61a���e��]�%=�ɱU����?!��Z_N.P6~=�u��^�o�X�U��%����M�k~�/K��@����r�S�+�����g�v.�z?bQ���q��u�f���b��a�����ݽ��xi�n��Z4�Rmw��.���X��o�ˢ�kM~�_�9+����o;%i�f�Gx���x����*��酢��	b�v�s��k�[���9uگ�v�[���&"��}>�+�?��bV�cE��ψ8��ao�D�szl�V�T�:�k��o-%Ġ�1I��rc�����آ��bKaM�Ye�R\�kM��u9��1+6������p����~ar�b��U3�=�~�䓬�esΝ��{{w����T�Ǧϰ�}EJ�b���'�[Q�σ[ҵ��M�4�l��߶9��	֪6�p�x/.3g� ���_2k߸��o�k;A��P�C;+����KOn���'/���mcN�T���4��t���!'L�L��6�R>�E*w��s%�|�7��[v���{J��_{�XX,����f6]��G��o���Y�m��5i�D��LG�i�&6	`X�	�B.����]��y���)�xz��ܶ־���rͬ�7w�M�'f|�Bz&ȹ�(F��¾�)6������E�ej�J�����g�������;b}a B��:��\���?�ɼK�&XoBj�g���C��]P���H�G����ǁK6U$�\�
	/�����3���a|m��B�Z�]��:����c&&�X�+��NOd澇.t?�u�R�<����j)PH�Tϲ�$��a��t��<��� ˿�d�� $ZM J(*[�
�9H�Ge���@J�M�Fm�X}k��=x��k�����F�'�cg
�1yR
�����"W6qg�� ��a��.�T1s2x�����A;�'��h�C��ɬԴm�*�B� �2C;��ѶL]�Ƿ�!����X��C����d->~G1�F���/�@�����}�Ot�����dj�1:��@�4�X���Չ��{bJR�D=�	��Ʊs�C�+��׵d~���<u@\ө�q:��s�xn�0���^g bs��}�d)�,X�t}����o0�����k1�W��k�[�6��0�V|^����7��2�����l�_�F�]�/0B<Zǜ�S�/ �!��5�`q����o#m��c���-^�j�r��-3<� �����U��88��r����ڱ�m�n���ffOA{�Ԅ���p�>������@p�S�X�T�&�*	�vZ�&&ވ�3y�4<���[f�eW��������&����^����X����d��;ʰ�� ;ݠ���� ��c�����;���rL_�G����6& p��:S�d�_��<��e�MH�~<f6~Q`����f'�ʳ��Cý
����4e��aT�v��*i�p���NB��ޠ��@N����h)�!s5�:�1���*o��i�%���uS��W`ʨՊ������j�G ��sF�I����we�$��d�!�Z4�G �=��HB�+\<�진f�Ob�����y�@\pMr��0ˢ*�#A\�#�^�3�D<�pkY�b����PW|l�=� @e)�~���qG�;��m�'��p��_��ݧ�����gfwd�Ε")��yj/z�l�k�,ܕhň���=�5���C�2m_K"f�ըR�f\��<�C�Lb:u����I�q�������������@'O�/{+�᮸S�Z��F��u
�b���g��� ��r�Yq�[Mr�J�{^��7�h���]���C̬��V+'�ׇ���I�����m=����n|�#*���C�x���"�ȆU�����
O�v%����4�����M����f��t`*v,"B�Z��NF�̮Q+���i
��fH��rǫo�p1E�[���k�$ΫoY���Q��o���Dh94kR�s�~���K ��G��x�t����J�(}G	�?v
r�^�d�/�lа��`+�$��Q�U��xm�y	$,�H| �yz;@;p����^xI��a�_��^s�_�D�{X��^�1+�[��0PO�>�ep0�;�S�I�e�o���^vj\�RŬno��_p+=��aT�7i���ҩPt8�9h���`�FW�R��,0�9���wn �é�����-Ŏ��P�1�v�[����C��)^����:z�'�_�dH�V��l����^�K*��S�z`�ṙ��8�PQ��	�A`��3{<�(����������v���l��>U�����>L>�sG�.�{�4�V�z��V�;M�
|�§͸��r��K�/��o���M�ד�U��N�����po�_�����4���.���?mR�-^�fױ(����Bk��u>��D,���?�
bY]��F,z�Q⢎��B��D�F���q1�ΣM��+�\h���B����"�ܣ��X�q���oL�.Iܨŗ��ŻS|�7�!�(�g� ��)�I5�ڦ�O��H�X���Zq�u�qA�Q���0Z�
& ��q_j�J뗇�~�AI�a����IY'�"�5a����n�Ϥ������b��~��tCwȞ2�:��S��S��_i�i���@�Jߍ���Y!h��N�7������Y��
���$u+���@�w~W���AT��6S/c���l�"X�Y������R�^�������q�}��&����Uw!:~3���R��B�O*m�'�_�I�Y�Ib�_�T��F����X��@:���O�L�� T~�s�Sw�q1��b��YT��"ԃ��r*�s�)��n�5Cq+V�,����N@I?F<9�lҹ�����t����aJe�D]������|2Uo)sYO�A ��������� F�y�I�I��^"��Ľf���m1 ���q��S�%EUOZGZ��F�;�jkpωP�%`I�M<�	hjy����#ǉş�@m�}���쨊��/��>{�.�/&�7�Ԛ;o�$��� ��,E�T��k~� O`x��J}�f%�����;z�Ol(�j�t�2�|I�} �d4)4մ4�;Q�
I�3��9}'n:aXex]g�d�mNT�qx�����;/eV*�Y��� S���+�C:<�V���.@��Й����������8���W1a���q����_}~��`��>|�6��׎U���FGY�1O��h�VwT݇��ȅ^�b��o�d#Z���0�휳E+�� q� i�C��}���p7/<��]{�+3�F�ȼrG���s'������&��jAH{�߶�G�\2����0�3R|(�b��TsJ��5�Es�c��ir���r�:/�m�y�J�mS�jJ�|c���F�ޚ�xV���;)vE�f�8J�*o_��پ�s�1�)�[͍�DK8��<�*�H<y���W�c����<+�	��a��� 3J��S�(v;��)��I�rL�&�����U�)DT;�%C�%�7��j�����%��9����r�P�e��b+�j�����}x~�șH�&�AK�MP�u�N3tk��R3Y�Y��~��=3.��?c�$Un����������~c�A�qw����F�h*���.]�������z�;���|�P�P������I>]1ӣ���t]J�$K����ᓑ�%*��f�-k�f��H�0-�':Wlf��]+!��u4����ڻ>5�ae�����F�<�͜L��1�o�,��.;��S�~��3�<僦����@����Ly��w*�����Q)2"d�y>��4apG4:
��O���F�� )q�0�̄a,�,��ͦ<�?�A󉟑Dp������oĸ�gLA�>Ȥ�Fl�X���{{J���^��afe��]�	j��l��E��>E����h�ڠ"S��u!���s�*��*��LZ4S��O���݃F�pp�:R��B�E�{�*L|�lQ�}:S��0�{ǂ1����$ XF���ђ$��`�e,ś�Q-�b�bn���S�cFDʼ��ĐE�	��x��wX7`|�����~������Y���Y���i?'����K*O�澕~8᢮��h_�I�h��8>y����e�a��q�.���%ts䅚�VִTb.����v�e�(PbL���^+���[��s4j~N���)����Uś�����x�F�������o'�������[��|%��N4c!������p�0.��ɳT5� �Tb���Ý�'^�A	!Oq����S���鏓V�
܀s���V��D8�P��-�}�����\Չ|�O	P7�g^�_}�a����,��w�E���i��"ˋ����/*�����$���L鄅���#��nm��b�yIb���L��E�������Spmƻ.����5�$��Rb��iA��c������
�Qtw��ʇ���RP��@q�	K_����K�յ�b��H�S솖�̀���N�=:�0D?�.���(V廜����ʁ�a'�j=�1\�j�$�@�l�Q�ݙغ9�lh���l�U�V-�����9���w����/�3���ܰ�!�O	i��a�HE��_��u�#�-E=�����D+���e|�Fw���R�,� C)͡|�X�ǹ��V�zʂ�`����D�퓦:�+hӬ1�����?��E��K͌�W��R�@1�R� �{k��ܼ� �KS-�����Ȥĉ��uZ��1�1�E�
$-�]����ϥ��V�	��1�V��{�JU\��ˑSM��9?�lsw:���6�Z�%�W���	���q�Po=L��ݼw������\']Wq��/��@�%��\�3F�l���$��pHQD���m#��Z;L�n���}/o�}؋�8�ˡ!I��l0�DSuv�\Ϯ�Q(��/���*:��]?B��|���	x|�ꉋ�)���-�|噍�f	�����T�E=�Y���;���3|�v����õ:�R�]7)��y�k�F���1�@K3{%��'2+�0�����~鏏�=�,�&�qkm�Xy���*�r��w$Y�3�������J��]�zFX��?i����a8�X7}yg��ϐ�%L[Yͧ��ˠ@L(1�]R8�}����P8֋��<�7K�����B=	���{��!�ԾD	�ɼǖ����LB2J2���ƻ��:�'�6�;�@-�ncw��♩D� Ӑsʪ��R�:�bCT�Rӛl^��X?��O�U�7�+�x��Y�Î����=S���:�'L���� e��=D�T����s�XT�c2]�]������@V۲͸`�o�U�&�eOy_�D��J"�	4�YaB/�ހ����0el���x�#@���԰�ЃfZv�LS�}�p�	���@ؗ���"t��� �;3Pu{�F#���;��1>���X��@P>N�"��ў�8��&�3�Ej�^�q/��v�پ�gED3�3c%��� p���7Z���o:��	M�m�单��p6ٗ�m������Ð\F�F�-U<e�	�L�{������1����M��;�II� s@����W�g�f��@����'6����qǹ-^}������(q�	�j�P}���̥M�� a�����[ݰ�6�i�ڢ�ƍ~��|�H�޻?�m����.x�Cѵ!og��;]�,
�]���My��Pd���#��Xz��/F��
/�֕��B����^�bcK���&����M�5�4ԩ�*T	��ʼ5no�R^��Z�.��|R��%<^�`>��]U�����P�8�e0J�٦s%��{�t�\��f��J��8��d$*Yu�8��I�%�����6���=X�o
��{�
H���*���)~"&������+z��61�&S(��N�k�b2�k�����
=�*����\̓�v��>�X�y��WrK�f����{��Qq� >��{m�⸆�(�_��ɪ��M�$�aDi£��7<�IZ/��;��\������IAc���L����0ӹ}H�]������|~�Q�M���n�s�y5��N�U�HV��yW�Y�#ݼ��FZ�Q�a�bGd�un���,���I;�X�����0C�&��O���<-E��V�$��
�j�"D�Z�X{,i3��7MS2����C'L����"��Jj�q��8���)*���e�BQ���+s`�/�X2��S*�s����d5nO�-j�Ck��f��$�lE�I��� ��b���S�zE1 _�:�V�����n��#�S6�"
��5)仴Hu�5�~�9���������X��9�+}!vXr,�n�!��N��!��en�����S�l��~��\W+b�?_q��+ܮB9z�X�k���W��I6�v����{��g��Չ���r6�wv���@aũ���8�>G��Ƴ�
��sGs�ѓɜ2�/��G_��E-�?]��4Q;©x	����1�7��80|�%ůg��tbk�?rp�\x={�3+.�Hf�b�4��Qv/{]&�MK�	��r cq(I�9�>��x�J�`!�+u�"�"&����
/�mKkZL42"e��e�,ģB����מ�v����Pߗr���+�~�е��I�w[g�����T3���L�	��<�o�����}gͳc&��R��Ϸw��Z-\���{	���Y�u26q\�^7bBg��E�O�V�)������p�΃����k{j��|�N*N/�+�%��ϓfח;��{m���D5p-�EB�L�j��.{��[�4�M�l܁meĀ}��"b����s�N_�/�_m����a*S�2K�q�/�����R��=�9$�l>9�P]K |-�+S��U4.�1�g�,��-df�]>&�%�{>�W��&Q}@1Y�"�p�S��S��/50P�q�j)�ٍq�w��p��ǚ�#��%�s½��.gҫ-�u�T2ř�窩�,h��ؗ�v�����d��+��}-B	��_-����d䌉��l����\�2�GD��_���Zo7LF�*U+��%3����@�Q~I�(�֤2,����[�����=�U�+k�֗��!Ƅ��"W���"��w�a���5����ӫ�>�b�x���E���>���@J�%���U��	S$��s����:^P']#�<e+�H(��3��Si��DE�Gdo%�����2"i�U3+���.b*��K�bˈ��x[�$�!��U�a�9�����O�V�A����@Zr�Y_���zY}�� pp*Qqm�5WdEO��j�H,�{���+�����u��&Vr��v��倭6j
����$=�,��P�s�7 <�Ѱ[ھStc������Ƀ2"J��9b9d�� 
��%�х�
S���۞Vآk�r�r�������0bt|ȗ?rZi#�_����!�7rW�LZ��ap0���#��=�h���qS&8�r���ۈ^��gOr�	=�g� ��٘�,mƚ�Ke����0g��b���V�4B'xl�-:�Ob%f>�C�+]ƅ��R�ˀ���~��i����v����.13��s��i
�����u�{�Օ��_F;F��4�5Ƚ�&YV�ѻ̕oґ��ں�ѯl�+���'�]�o8��`����f�M��$�٪q�o���C_k��-�o���u�W��R��\*߻�%��!����網�*�!w�]W�	��|(Q$�k��Ŋ��w���e��ŕ�	2đrAz�$.!8>�yN��q��>���]L�:�u^�������:Ԧj\A&�9ьɠu�
�-׮U�{�UG�*ꃶ�D�ĩ��Bެ9��<�2q7�qm�V~���m"�΅q竔	#���H�[z���'�?�
�~�����Vp���8��+�N����T� _v�4J7��qJ�"m�#�B�u�)Ĩ����]�>�^tL>H]I�m�Z�C��ί3��|H�@� ������LZiy4x�l���h�/`UV���.��>�%�ƗY��2�oܬN�o�(\������p���8׽.'�b85S7		�0�L(Fq;&�Ti���C�X��Lj�\�G|��
@�������$��&��������!W��W�q���CD������!���S؄�� �!oM�0��_�qBԑ*�0��+��q��7w���+I0Y���.#��|�KW>O(4���*��l��$`F
?~YP����X���4�t|�@Y&��h���3g��������[d]�ۄ��-�wsZ!�9����<�鬚�,�$�ۭ���8�O��l4ix%f�E�ۢ\0��p�p���
�H�ĺ��n6��D�W7E!�PBJ�����{Teg���K*_=��?t���5�<g_�L&r=m���=���r�On����͗S) iPW%3�#!���/� �z8�}��T�Hu
-��4<��?���o�$�O��U�2j:�)�Y���f�>��*p�)y�HPݮ���oF�|�n���es`�8�ʡw��sWy��a�؎�� �q�ƹ�`��
5D+F�Y6r�N7ui������ʛrxCx����u6u�`�Ii��z7�F?&s�7��Ӹ�n��`@;C��D+'/���K�'z�+5�����@�R�S!2+���v� "egD�ՀC�{No��^�y�	�Idf�hU^��z��S�H�8,1M�%ͯVbO^i�%C�O���2���|]Zo�r�ϱ��R^����M��3%�7p���JƎ�:P����mO����v`P���	���9F/=%�_n��~�䪡͊�1/-V�I����Z����gw��	���˔��P�s[y�S2zç�*�����X�j��9��ӌ�jI��(g^f��>�/�|1ė�{�����7����O����T�d=�=�w��ã+�]$lZ���2����2��g_�BȉE3���{wt!D����d��������.l�!^�s��u�9�b4z�kmZv� �w�- ��6>��;<�`�VDX�|ΌX��|AoJ}V��T�X��ۧ����)��C4��!�;�C���h��j=�44<LU$>�8�O�ܛkBC�|oy,�s_�G״������K��!��]�8,��	 ������]ߒ�y��W5S;Us�̱���9ݽL*F8u
R�c�.H.�h���Y`��=2"���W�,hh�������Z ��BM�-�q���ԡ��<�������ۋ�ݬ`R�o�`���7X�4ނ*�S�`��R;cQ�mB���H��h�{-y�y� 3����jB�]07�)60����%m/BхСTc�ԛ��6�:$�g�|[�Bn�R耠H���:��88�?��i�!�c�ޞ�B�?Z��Ю�A��6X�nˡ,��6�_����&q��󰊂���!��}yC�=F��.-i�#˩��|4G�����0��yRi�?t&妇��:x%O��q&t�i���u�I��i��*T�4��z.7K.�	����Va"�lj�Aɢ0���� bH�Z��h��f5~of~��8�@C���!�N�J�n��Ӻ�w�.~�v��5/���.:�Ա1�Z�+ڠ�?`S�� �v�Cݗ��E:��,�mt-m�R�y"K*���������l�'42����![���T��*�.&�Z����J����������w��b�?���m/m��q��@Y��+��n���'��e'��<��nW�K�Xc�CK��S��}B���.[>�q��gFk�W��#�!#1�ٚC��q�>�;ҽ�Y�ج�E�����2k.>=H��2
vb��*�>7�%��2�	��2@o��fG��7�//%�yGW
r�jW���~T��Jnxoxd0�A�(_�,���ݧ�j����z�ؾEA������h�][��w4 ��}�,��mM���no����ͺ�� ���ď���c�cK�L�w;�ʆ�A�՟���vSʄ8�Z��s��w�]��>.>;b��U��v��n`��-�zac/QJ�|�1��E>Ԗeu��%���=�."Jun=,U���[B��U繺�έ}\��_�l��n�d�u�(�8�5aپ^�ͤ�W8�e�Ü5�G����$'R��Ow��u>��ñ�z��ng��k�g��<�T���}HWpu�wJ$���:q��tBe�]v�9W� У�}-l���Gcُ ��H�������[���9�X亝�����u��V�Zy�
��	P�^�l��RB:�BuF�� ᕆ�H����~����ʞ��p�-Q��M��'H�)���d.�s~���?�R`���>���Q�@o��x�`E}P�.�iu�ab�+&3������݄z㢪��qX�F��!��Q��;��4�O��Tߙ�M���=r�O��)l���~� �.s/�?��ݓ��G���r��x�7��`�شc�_�M�i%�d˄i��:\2s�� $��sڎη����B�����<��I�����W�/����v��6����.1�:'N�1�Vڷ!�o�b��͆5���� a<E��S0[�&x~P5V��Q��غ�zO�zN�TE�qcVݯca���f�Zb�(�)�a��&�]���V1lVg)�W����V����aVcT�5U�ֺ��6�E�F�F���2E�HJ��IWx
3aT���ڞ�fvQS����3/����u<kH�x,��e׮�x�T$��Fu�j��Q�lȘoW��R�%�s��`�VyH�>%M���I�WD`ty��]E k*G��%q׼e��T���Shw����av�8�>h۽R=��^��H�~�2�B�b��a˽�?ˍ?k����@�O��\�m"�p�oz����=)4(L}���[�5�gmm�h�Ehr���l��> �M�s�����h���d��!����I�P���f�B4)g_s�����H7!��E]�b�O8<?3xM��]_<3���	#����h�,Nk6]5'0�MzU�����/'����},�˧��O�D1Vw��͵�G��8��)#�Ѳ; �5�� ���^�'����"��%�o~&��լ��yyEmA#e*�1��h����|�B�{`eM�J*Y/F���tis~*_
�J�~�l&���=��Q̂��
�[����Q�u�(cL�{'���$�wġ���n�.� �2�pZ	��Y�P�r����N����-�*�\��d�/q��om(��F��J��/�Nz�=�-YtT4��?L�`&Ҙ1Z�o�N�n��:dr�������2�)���5�&f�N�2�� �*e`c)���AY'����A��Nt�R-�_{	i����X6_��G����,`�3�[�c?��SF�}�Sà@���&���PF"g����޳�ͺc# V�ި.�?m���8�ڦFed8>'H�]�]^��D%ㄏ.��բ�rK�|�`�g��e��9r��ӑ��2��C.��XS���Bb)�f&����8L$4�$B��O��S������s$6��N+%k
m�+/����:Ӱ�*- Ã�x�q�pZ�4q*��;�M���ۭlTCL��D'�r�7�9<3�}O�C���ዖ�9O��:]�k	�Vj���m��� &'��wsW�"���Z��R�.����]����ިU7_S��l5��7Z�'ⓛ�!���}���C��?�Iz��?v �#l���beܐ��p���)hoO!�l��7л��E2c��w��=عe�
���=�C�`�s��dl��=�ҷ0Pt�^b��>�"f|u�69�Ÿ}�(l���?��K������HN��;��[�׊�Q����yB}���ˍ/�;t+��4��|L6o%���,���S\��v�!��I���Ēb.ø!��*�O�ڹ�E5���-.[ٌ��ܼ���蜮?�]�>�5�(��EY��X�l%���x|6�X�c���|���T&�0M}@����7��6�R.���6u$UZ��d�7Ok!�w��2��5��E�##m�Z� ���FkK y�]O7���E�Ո�@�B��:�]tR�@]�6�"҃C���$����`-��yj�ɿm����~ݛ��������hi�a�2�T_�^��Y�������䯂t�顷AA5I[�mb����� ����� �	~��'z�X-̺�n���N-)ٚ/�A�s�������?��q6tp����($t�ǲ��&���eN!P�6�M���xO@�8�$qd�����`h�o
LڜϮD��3+�b�����w;�f���3���ċdݢ��R?��K>�&nG���b�*l��Yi���Zj�龾p8�����7��I|�����*��J)/�B�F_��{��2M��v}�H�@�
�iir�<��h�<��AT�K�x�-g:z���Rtx"�5��
~>�vnco_�5&����xDs/��$h���F\�΅y������5!�6X6�>5�(
�/����u��҉	E���~�rB>"!���E9����G+L�f�KDII�Ҝ�g��q�o0��*?u=翆�H��[��V?�I��s��u���?Rq��&�J)��H���T�-�8.eo]t7���9|sbb�L)�����'�N|�e�M����؎����K��D�a��<m�L|�)瘈!�+_U=�@�QѴ�"P��q�;u-{�_�u���m��h�[��eR������U��a��L�u�p�/3I��3le��RFZ��rR�4q7�c?���w�8T�˵L�~�@�������5l>�&]��|U�-k�ou�On]%Dm�c#�^�u�>�4��i�p�����Z�#�]���$_`h�J�ց�_�q|a���������p�<�<H��eC]��xdW.�3G9�èŌK��8eO��>i%�+��q��Ѳ*��8��9��%���`���{Qݙ��f\�T����1^���>m��h=�J����b�y ��s3�į���>���αw�q�d�)��-|�A�d�e=s���SZb������Mt_�H� 1j�{�����յ�Н�Я`qMD�}+����d�d�^1�@����������|�q�u����V�S䨼�;��&�,��?~4Q��_g�q@y&zb�L�Y�<���g���#GuE��������i�	�*S�����٨)(�wz��'nB'w]�n��$��5��	�0��‍0��O�����1s�?-P�>�.E��E�XqNL�=�'/㍵�qW�qt���Q����a�������$�3�4�ټu)����b%l�K�+V޾�&�g�6n]ַ�ӳ�1��U�����qE���?���������@��(����u����2�'cvZ9�/�R7���*�f���"JI�����#>];�/�>�o���^q�)D�J����mO��/K?�^�i��4"���d����u�Ҡ���--�NE����[Y�,��{a5��V?�p��]�eV�������M=�o�L0����+~�O�z�5Y���\��"�������ֶ���3_�g��qi<���gC�v�s�$�qM���3�T���R)��J&��w	�G�`�7����R<��N��ݤ#;ɪ�&��j<lB���Ƚ�	H��y��|"�t�qh8NHA}#ϙ�Z/Q5�{6Y��Aިǫ7Y�l�H��:��d����K
I� s}+w�4#���"��c�*>>�G��}n��`���"��A��B:���PO�H��)��M0� cQm��X�v���5�N���Ȝ��H!k�2�vr�A��ϊ�?�\~�ow���W�pD:�}��p���u=ꍇ�h���TAA�$��P}oR�յ���^�,�����
`��������s�Ը����ټ��!M�}q�����[xAG�Z���s �V�/�˗�?{�}s�'fOSTm�%���jeJ���
p����	N,�����ʛSaХӉ�@D���(���SE�{�R�˹��7cb;�`.�_��Eڕ��B�����ҽV�{���Zw-��;��Ƶ�F�v�ݟ&|��֕��(T�J(�&,B�d2�H���eJ���6PR��1���^���H��Mt9R馀�G�WqұS����yr�Y�@�x�c�G�<�+� �P\T���7G����B��<qC��}�~ۍ-$����_;�\��Y��>�J!�B��h�ge��Tj��o����+ϒ���K���sOA�M��b�߇� �i��x�
�	����X��
3NA��XC�"�ˊl�z��W>�@����J�R�`��㟁��z��T<ҷ@��v�bM#�s�	^q�FA�ߘ?x����6���ո�͢�1<�d���|���'z�ۤ++�����~������� (�+�r�~�T:�X�tc�R��ݫ`M�]�ao�-ɵ�)�&jO�W`�֞�!0��v�(��kWCJ���M�����W��f�Y�uw�R�5��нs�^�Q�{�X^-y��1c$�?�ר�E�a!$0��q�Y���A=.�����G2*��5���ټr�D{|=h��v"�&��_g{��׏x��jF`��>c��8�ς�d�{���_oC���u�U���s�`!^Ǣ�b�������r�P�컑�߶�&cG綥hyT�m`\+�_����kj����Gb�䭭=RAj�h�?u���	������s�:Y��\J9�n�L��q2����Ao����_��}�����Z�)�iU���` a�����_�S��k�^ƪ�Jf>��6yN=��5l�@{w���Bli���3�q$Ė�	壡��k��x�����e~�~�Wji.r��`��f5V��O�� OO��Fw�~�P��'6T�5`C���x������~�*0va�౛bjL`) rXJ�T�ᬬ�=X��0Y��R��b��B�c�h8�35���w~H���<"���2,�����LQs��W/s����� Q��¼�"�y	Jh'�:�}F@���)�}ʫ���Z���-X5�vm	+��"k��eVO��w`�'M���栁����|�X{�o�t�0g*ѵ�����/ �M�V��@�T3ʱ"W�N/d`N}��)S�K�{��E����e
����Xg,P'e�#���u��K�$�,뫤�?�����D�Z���|�|D+�,K׻F�%�Q�.+C�8��	�#�+8݈�v�P2x��~t��"�đ,릣:E2���)H�1�"`#Ĺ�U�u!��}��=�,;B��H���?͘�Ș�x�D@޹��k��G�c�۸V_��d��`p>��sX�����eLK/�kˑ1;�Lۯn��:g^-�����ﱦ8��F�4���\ �����?w�D6�w_\�1�pk��K~��'��t_��\&X�n�:	�x�b5�b�~�Fx�V6a҉���������d�� ?�FvU��x+d���H�f���&�_g��/v
���TkX��[F�z��!iu�}�*f"���6��{~���ȓQƧ4���a|!�o�E]2U�+.����+W�|��/�٥�yi�1�>��ނ�$�?�ῄY�G� �Gb�����6G%\�ޔ�k�OX�[�m}��p{�+I�����"�^'$;xl��%a�h�#0�X�I|�/��]�G��A١��(Q���-eEBm8�-��|o����2@��|�.�ɠ������T,h�18#��\�9Az�x�N�4�Ě�[�;2����}b<x� /��^���i�M�>��2�ȶ����6�)�e���ɯΝ=N��%��{���Z���NT�d��6������@�z�E'Wo�ъ�A��3�y�a��	�E�Of�Ѐ��� �����Ȅ�ٸ�P��^Gb�$��Yj�W�ҷ؅j����k��U��د�g��3C��G�A(�~9�^��Z�6����I���o�)>[��3�gr4c�@��je[�;�©���?�ى���p��IR3z�-{���R}�ۻ��م���vfMg�z��ގyP�os޺��o����?i�F��|v� �E�@w=y���zR1�S��t�J�6�0=%]`�N�;a�0J�c�+�����=)�?őw�I�>���0����$���Y����r�-�i(��{^mla��я��o^n>����&�U�`��h��ݶl��*݇lj%�(f�����#B�ѡ�d 澿}���S���6k�r��=�v�L�	 <+�M���J�m�:��FO�u-�II�߿��voc��MY�O����cIN1�t��0���I�\@gό;��O����c
�����1�D�J�Z�
�H1���_[��W8w\)&|ϳV������}<���.LP����=�Czc�`L]ب���%U��r���~Z� ��qC�]	Ɏ�>8⻞�[�"���-���F��x���	B'���e�am>1r:���k#���?�'�q��o(��q��w��^O��$��~Π�Y�72�d� ��`�=��U��γ!�N�E�N�F9�����"p�޼�(�C������e�؂Di�l>�xi�A� �.w~�z�`bG��OD���r��{�`x]��{�4Q@�sJ���΂���Xq,T���1�FĬf�o$�Ԩ�>FI�o�n���Ƈ�.�τ]�����ƌ&��]�E�iu�c)�ij�N�oJ.*$�EK��ju��e|�ؒ{��'��~��������co�p7�A�XA���������Ĵ��s�G+�/mth��g�w
>���I��>��)��J��wbqb9�")1�K�R����2>`��H �l&�h�u�(��R�B�P�4��@/�Z���AS1۝�?LPU���*4�b��wQ��y{C.�oc�-��dH<[�rP��hF���F?��	X�9*��>�RP:f�e�z�T�Mn�����#ҥ������T��f��}���oAt��qף�@bb_��$Օ�	Ĳz�u�&`ėח��7�D6��!�����W���oo����_=�ll]�F��m��ӆx8��^�����v�UQ�� ���I�_���	��U,���K)¿��m��2��5��y��@ܽZ��F�:"��s
%n�NQ]���\��2�X� X����ý��n�K��f4щƿ�f��U�����Ņ�iLN3��i����ڏl�r���	�h�[x^cH��JL��^�h�����t�d2�nJ!��TwK*t�7�����9Z!�P(�Zǲ˦A���3�W��s�i
w��5�N�ǟg�� c�Q5ǂj���KmgΓ�_~��9�����#m�[�%� ���G`b�u�����/XҜsޮ��b��+�xB&��B��J��C�2kٲG/G�&���q�4�`q^\d80�wA� 7�0Wۉm��N�g��oA&v��?[a=~:���Y���L?hY�T�V�'Ö�T��W�"�۲J�@J�IRd-��u�Z������$�PIT(����HV,A �ܩ�Q)�2�!�J#��Tڟ`��Quxh �(��LO�s)݋�?�OA>��۴�K��0��b�T�Ϲ"hM�(�q����O��pXC��A@�3�y�/���_�{���S��I�ZA�O
����"@z@��SS;��&G���'�U��*z"y�_V�X��ڌ+��T���k%9ϓ)8(4��S	��5&�� �N2��?��?0�8K��g}��,��HM�M���P<�쮵�zG����vG������64�!�.ۓyr�r���Z�W�P��?����7�Q`�/p����%��S��+���+�?��$��#|�򯰜$��������t��V�i�е�$_=X�^���S�D�L��H׎K��Տ����;b;���^� ��>�_��~z���!2�̝���G/�y��:|� �Gw[��<�M��h�4��Y����,c_���YȮ+�ꌢ����L�l 믬'�����Nr
�֍��k4?/���P�dhw?uj}Y��M��"�_�r?Ee.N��L�=?T�^��v�r#��8��=�=~$�a��S61�et�$O��_r���y]�ڀy��o����ﰩS�/|��Ĩ��Z]v���}-=�a�t
�5ձ���ԵxY�vl��.�_�����[4�V0f��v�8��֟����/'#�~L���Tf�G�{�ec�!P8�Q�����Y���B��O��,pE�����"�N壊6��65�$6{�~�2�l���c>�4^��(¢�_��+����ާ!\�d(�u�Yʃ��Ť�r%&P���� �zȰ?��َ\�uϴ﷝�� EsJlQ˷���/o��5'����P��6=��2ZrT��>�8Y��x� Ɠ_��e&�'�/2����,d����̝d`5����a��n)�ї��-��،g��P���k.+(P���?5qn�~�dc�N�].Gc�c����T�L�������%�\��
�T6m����arC9��\:P��.z{��s�tp �����	
u�ϵ����d8�� ?�K��b����9�w�]
�
�8��'7�a��C(L��8��,�u����f �T�9m�]?;d�F�&�4'��cf�_$)N��-��d���l#jat~�j.�JןM\�~�����/��1�� ��b3�8�T$a|)s��:쇅�DD�Xb���?���L4sAh�*?�����>Pm&\�����ϐf:VM�G��22T��rը@�M A*պҝԕ�6;�'��+��T Z2���-Ѓ_�Z���������K�M+�Q����C!Z�؝���Č�Y?�����h�Uk:����S�`T��G��yl�4^�X�?޻v��7�F���i�����${�K�,�m��,�#t�����s% ���W���C�O���HJ��B���q�����$�~�,g�,a8���-P'��F���Fd�W"��4+�r��/��%���� ����BWh
w#�BJ ���􂣭�͟��:��.�X�#��>-���?�=w���)\�͒x~tڂ1�'&�䖠2��U]bհ���c�+�M�q� N`�:WVRϪ��w����8N��2nd`R�E�,Y;�e^�&%F	5{��'S�J(���S~E�-K�c3w��I�g]*`���"�o֧��kO���5:�$#����	�a�"׏"����ͦ�O�� �Y4(�oPi,�W��.A������-S�k���g,)G 1_x��~3���� `���7��a5�����F��,�	�ˤn-�j�TO�
_�S=�G��$��N�F�A{�h�<��<��<q��F����\(o���ܸ�d��&W��uE���?V(T4 �vJ�=�?�=���@�&���|9��5J8*-2#m4���e���9��r�6���C`@g�OG-t'K��l��E����]0� ��4M�c�W���y�J08�2s#<�3|@���8�>�vF[�0׽[uh�NX�p��_�I�d�U@���W8��x���d�#��Y�S�p��-NQkh|)�U�MJ�J�RR��k `��"�^����㲲8B����JB���BL��m�X��o�B�!�ϑz����1�!M������͗%���Xur���-�:��J��|�]�u�T��b8}��}Z�7��߲��Ĵya��T��_�̘8��ӎLÅ�!�S��*�?���}ǳV�Q���~�P��K:W�b���o������j�ځ[Mq��-ݝ��8��S���+�U{g�Qr��v���r�N��zsw�[��yid�\�.�X��S�L;��'˘LQY���{r� ������,�LJ�	x3�0]R%iX ږ��Y]�%λ�8{̍��)�E��*�����Ч���+�K�m
DZ�-D��䬅w���|ӎ��8�b�0.�,�~1Ȥ.%e�A]��e���
��%�Ai7�g$XU��s+��~�( 9Ѹ�嵔;��� �Jm��j��J�MH��*ч��%^s�F	��8
���Gen�܍�l#I-JHy�Ⱦo'�J�'<���h�����rNj,-��{��A�do��L=��bT�?�Y��FO0��������~͐�<a9����6��oTPǚ�%�V�h0	p�� �
�1ʉ��ƶ�x"o`C�|��Zs�'6W���D~�ެo�NfD��X���_�0�w�ظ��V���{U8i
�ٗ��idn��xG�2{_��,��A�:c�Rx"wo5S�E��k&��.]�����f:,WG���4�A����)�꽣и,ݐ� ���G���(u������������F�����I�!E��{3=T�>���X�9K�b-w��Z��b?L�)�׀�KI��>Hkph�7��DSl��u1��nv�z�����$�;E8��f0㚌	၈VB��z�0	0^�RZ�_>B&���5y8M���Àl���&$F �� ��}1�Dx�&�Y�P~��P�L�#Q�������;�}�4��>�;�~���&Mwe�ܐ�ˏ52��U�D�@�;�u�'F_U��Xq샗Bt�3X;�Yݖ`:� 0��~��	��0�q`�V�����BŚ�3�+�F��H*L[_Pu�}?79�~��lo�xL+�q}�L�P7��A���\����sl���T��jv�����V��C��{���|O��*�y|f�V�������\6�z��j�1q�V����K��x�˚� �frQ��.7|�éoP��Nv�^��o:/	Rp'��w���".�DV��J�5r����/,��(ܢ'� �ۍ�ּ�0�Y�߄y��#uR`#g���G�~W����p�e��Â����J�GM/��A�P��^�l%Y@����i3/L��ݼ7�R����z����<R,}]3��K1xF1\I��Be�~�+͔��j@=+�Ϳ:���g��-��c>�t��~]U]�؄��9���/���vt�_��M���i.D͊d����T��7ܖ����<����
W�����s��As2Y ��vOQ=��m�>�)u�����u���+�mw�:0��sR�����n���V.�A��r&P����4�8Ws��o��3s�Q5�n�@X�:J�ac^������~�@� �j��`Y��'���__4ʠ6�[]���z-%wD��1XI����|}�HҬ �,�=\|Ǽ|����J-���,	��B�����_�@U���3�'"�$�,F�`�)7��1Q����$�����������}�"β�E�V�@�u��-Yф��q�mk $5$�1�H2���}Ԥ�I�$x�pq�2Bt/J�^�j\����S Xj�M��g$�G
U4@�S� �>��%�������g����� ���T[�lD�j��Su��~���P���Pq����9=�uIFqj"��mk��T׌;�1��	ٞ:�f��Z ;����B�a/V#���yZИ�=��\3���3�5�J�)H��^Y)��wLg~�T���(>||G�hʼ!l�H�d��1<����G�����~���X\1h��	�FV��CiF���dD�ђ�D7��(�H�����X����E��CY�ċ�QMi�0��:���	C�|.��ap��vj��t~���Ph�l"�.k�E|��4�k����_�`�� մ�wd�Eg�#r�e���d��<��dֵ�����ǲ@�jP������x���^�QF4��*��k"��~Mh֏j,˴e����
�-��?u.c .r$�Y���_IL3l2��r?����-��
�u`c8¤,� trW�\6�²�]R�\hf4;�"�.�1�����*����s���ІM���\�@��{N?��	�n�~����������������}(M��rj�h���[US[U�H��I�b�(h�mM�WN�	��ɜPC��94}g"}�Q��#v�ߟ�
�����8ߍh�}E1@��(��J�'
W��t(����v��R��<^ûG*���2�n��{�6�g&Nr���A
�D<��?��^xBp#� �Ҝ�a`�����2DTl������������j5��xq�ؼ�̷-�|d#�'�W���pw7�Q��j]8��y�HxR����o��վ�,���QUSN�0l3Q��']�ٴ�S��O����^5�W���t:7�fĨw<i��<4I�d��S�������"�bp)X�S
9a-m�C:�l��r@|�F��㫑�c���i:ib~r���n����3Y��&�Cʓ�-��7P�x�2o��31�U����\-��m`���'���	�:��#u�
��q	ń����$T�ЇN�~7b+���������V�f��CD����(��Nk;�U�KQº �����4�9�&�M��M#���_�i�����Y��qƳ�`*�w~ ��`�aBU
��=Mqk�A��`E���oM�J��GKO�fFj�&wb+Պ	Y
T&�Ƈ�=�D��[)�	7ad/��R�7�����i�m3����쳽P��R#���tC�@v��w�	�^�TX�V�H6�OV>G���͋�@7�5�U��EZOխ{��Y�Hek���0:{�p��&�_^ �鐸���>��$&KjG|X-��@�>h�[�����M x\0S���1X���vV��� �V'�����6�![�h$ ������V��r�/���~`�G�p{{^2��Y�:!Kr}��	��5�7J�e1�q��>����`��|좡8��jp�QQ^^���#��?� �����_��;�ԙ?��.T�2����B�$����\�}������q��FT<w�ɎU>f���%�f�)m�i9��vk3��eti�FE0šLbY��o��*#,�t�`K�����w�E�(�0>����9}W\����� ��P�"C��c\f�'Q�v�������BBWC:�6�>�{��͠�Þ�Wj1�G�q�鮓ݯC+�im� �Q �ZD��:���u~��عA_��$���myg]`l꧑`	F��VAz�����5���M1��9r�F�貃��.Ã9YB�IT
�]�:�?Yk��):=x�[�$k�@�-������0�z�e$U��mz�uFOZ.����L��цH�c�ľ�!����DxB�2��[1��`��>'�[�h�Ǚ�ȗ`���3�~��Z��W��6������̘��H�H����:�8-M�j/H���]��;n3�!�q?�>�Z͋���������MP/P�p�񬿧J8���G��X�q�����@�Ӌ���g{�Ȁ�.4}�X�5'#�{'�c�F����t=Ʈ�Vŕ��9�<h�?���IZ4S�ƀ�]�g��m9�&���9d|��R�+�Q�������WG1�41s�[o���j�*z��WD��
Ǹ!�	�<�������Г10@��Ƣ ��8��Zl���X�O#�V2����ψ�)f�h�2X����q,��ѱ���B����hWR�i�9��]������3��ױ$9(Չ)Zl�E���p���p���0a��&��S��o��!&���H��#=�6d�ypc-;F�W����I�I|+E�K��I�m-J|0|rW8��7'*S�>i�J9?��/o��B5�U�z����1��+tq��|M�T}{��b�"�*|^8�:���c�����O�JE�U܀�0�t}.�K�#�,��Ä��v�z���e�-^'z[��b+���N3�X��l�>;�EKK�GV�'�|Vq����(��َW��:�P��v$��,ҫ��mz�|�:U�4ZY6d��̫�d��G���2F&x폧����"��{������=l���vVoWO�Di�ÿU.�g�/�Jaȴ9s�4�!� ��y���A�zYy�0RRl��X�p9�|_h�J��E�&�ǧ��eRu��EK�TT�t<�=��(:j�Dq'N�#`�< ����4�n�j�R��E'Y��^�
:�y��{�����$&'p�+��O��X:���H�a�\3�;x�w�,|1��\��Hr��qA��������v��*��e�$j4ï���}���b�>����^n�"�����F�<t=����шQ��������.���=]���`��=�PP��W��(Ğ�]r���en��Q l���̵�����3G����w��Rq9�K�����}�UAxg?���a?�U!��k��<�A�S�?*� /-�:k�G�� 8&"&K���۾�˞;���"�/;��m�!��?tT2��y���*��`I��߅6@C�v��X�ڭ]�Ş�|�,��L�Ҿ����m]'ŝ�B�ͧ)����5~�|��{�1�{��!���u��ʽ�jr�U[�����l�,rE�v���r��gѨ���	�vkcW���~T�fz�hN-�m�7�Q)*0q�w'�`Q(���\3@�J�-[�僽lNM��4b�ߍ�#W��vf �1��q����G��uO\V ��5u�����6v�ǰ�W��l���W�t@��24m���-cS+qh��kܾ��ŋ�����	L�^�~B�.�b �5)�帑�>�>,���MK��C��|#��,V�A@%~Q/�3�׃A�\A-Y�?Z��R�,f�{��@��0>Y*�w�CŅ���1�T���U��������F0Ta��q��ʍ�o�����	�9R<���6��?��܄Gh4���0p+��������o?Y�A�T!�\�S�z�;ÕW*<�1l�����������Y��GS���~�<o�Q�0�R�f`/I~#����_�A�9�S=ROޯ��}s'ǱZ�ة��9Q�=�]i����O�E~��QK�i�W�-]��D�9Q���Ev��K .C�J����Z5�
C�%��x�(�����@����+g������ֿ�C�bB�z�+�a͟��18Ioa�a�{b�OJ��/_��)�p��x���q_���)�D���H�*�Fģ(��n��:��=H���u� �;�T����Mk�^&n��������	]���ع)�e���[�_;G��1W� +5�Q3}ڗ�r����XK��c�?DT���i���7nUoi�I�R�2���q�%	J�J�|��Tߐ�C�it�>V��dB�8�έ��y������S�L �.o2&^�(OG�v�(��eM��~�87ݿ�������5�i��2��n�g͑ ���;�ҁP��e��R��x����`�P�0�6Lt�-�Lt$�M���*,���ݦ�.�f9��\cƥ�{}]�ߜ�w:�u���Uڙ�R�8YY��M��v&:n�]���M�&��4��?p�Q��D�?��x�>�#}}Xo�mAN�1�#X��/j2�F�,�ʃO\��t��TJUe�u	���q���Pj��UOG�%�&�#?�*�]J�cWM/;e��.@�Á�gM����Y�N`95��	Wy�ܔ�:��	Y��&u�1y߃{J�'�2�O;4c��U�Ų�)p��B��驅���#��-�E��L3�M�{nñxQzz��˕��_����[`R`�� &U=1��S{�R�fc�9b_Ioo3�H�\�־��u�o��8��Jk&�;��L�-{R���<�[%;���?��9<���zc�q6j��6��m�vۘ��ƶm�jؠy7�������d��[�>g��Y��D���&R^��W� �B?R+l�Ð�w�u�a��Uֆ�X��f1���j�T� l�l���	��ʉ��4i��c�E��l+�)@�]V��r�.�.��3������:ibDtm*2ڷW�:�}��Q���lQe��Wy���˽��x�ώ���_4Q�(n�3���:���]�	W�|m_8v����"�I�>�;N�e� �V=��O}�=3X!���F�P�@MO;�@?�l���:�5y�Q%�ڏW���Oi�S�ZO��ɦ��R�ߨB y���j_+8�*�juLrj�5[�zԆ�퉵S0mޤ�Tj�C�vQ�\��������;�FŌlv��W��+%��t��_�������������W4�t8�-�L��P�!� X@�r {�2ב���v������yĘ����o���!]Z��~vD���F,��FN÷�$|��-�>$RZ�~��H�w�4fb��OD6'�Z�Zj?��@`�jk|��������8��f�{zNd�2�������E��{�ȁ_���Zč����~ =��/;uz��1�Ķ�9=V�I9���29Q�)7�J���7��2������ܨ�/��,�'�-��$k5 )4���?[h�=sk�yK��S��B?-��+R��wi��%��;��x���.��\�7,��Z*'ޟ�*o��,�1�2x� �W�4�:Hws_K�$��;����L��	��yK��v�S���չ���I��HZ�(�i��Ռ���W¾�_h/�#x���D��T�}�ǽs����苼~�>j���P�)���A�v��r���y�Jj�&5v<�0[ۍ����p�_����W�-m��9t���5>ˣ�"��X�;B������wE��w}ǽ�mŶv�8�4���f�6h�-��T����Z'�qJ7�,�s%3�S-@�wP��~~]�^�&e}�2<8X�;��	{AP	����/��=����Z�j�f����Oz�M���~s$@�~KA�Eψ�ɯ��`7��7�Y ��N�j����� 3���T����ᖻ�"|�x�DR�
�hr>��tG�DI�8d���	!u���+��Ȱ�8�U½)8A,}�W�Y����;h��5���aP�� ������+pYS���c��
���Mg]?��o<�����-�3���������T�V��k�+e��Ӎ�J���_�������ޔ�@)6�'ً����j��� 	�ɫ ����CN	��+�R$�.��7�{��������}F�׺����7�����u�����C�fZ��3*��Ʒ��*wO�Dw��v��
��� �8���i���J���]�{~ m��y�,���� �`2�O3`c�
�vsO���&�b^�=VmG��'��QǹߢQnS[Z��,��!M	��n;i��C�k��i_m�myG� J%K���w;��K7X��3я"���Z|�_(�x�M����3����uZ�v]�%��@�J�T"����,�!�,+����K���u/-*���t*��a%ޟ�J�[�v*r�G:/]bk��i���O�6zLiM�V�����t�4�mG!���Ԕ������_3-T'==;�Ϡ��%"��R��Ǹ��V�P��!��>�u�FS��bi�������}�k�y����u�z��yv�y�F��+j5tn[�2��Ea�n�,������3<N:Z�O8�\��z��_��KL��9/C8�/OCt�|H���t�)0k�e��r
\��_��?Ԗ؟���*�,�A�nz���y��� £�ص8��{Z\�����-�(���ӿ����d�Z���7����j��f,^`ÇL�u�2g!"����n��� v�^g�)cN�R3�V��C�/G��>!�A��A�z��+��1���ȿ��,a��CEC�^po����3�~��c�+�[�.�������͐H�u�ߘ~��X�#�
��Q�� ꭭����%D廧�r�7mSg����J�����A�t4���˂����^��Q�J����ӓ����;���fBٛ~��I֛��"�E=6X��~������m���;�Nk:�bt�[!{눛�T�R�����`9�h���,B�̻��|ғ]��;�/+���=R�cI�x�o� ����a+f%t@�;U���/�S�WTo�L����(����ٹ���N���[9˯�}������R!�?ɩ7�����-��{/�z\�/K�|��X��}	��eT���{搑�P������E�9u��]w�r7,C�Eqn�PLj���Gh�����x���Q��BxUVZ?�3���_\�ϭ!rT��'!���ż�������rY��у+��7��iyx�T3#�ӗ�o	��󰍜،�H��J�p2�W�/���P�x���ޏ(/M ��O��R���z9�� u�~���u�>������AK-p)n��-����t����6��sj������.:���*<�r�B���@V3�����4<���㺪����ʒ��m�H����O�	��u�� j?�J�|Y����`�l{{,��	<�U�!�&���RWKI�;���<�6����x�ʹ̎�ڂRK~f���;��s�a-d�y|3ל1�S���{�^�z0WΔm|\h�г��p���!��Wpat�P�ӭ�����~�][$������Hf�]�θ�M�-�}�Cw�J��e�;Uk��j�e(�
#�����Fm̧@c����=|�5ՙ�X��n�^���Zs:�W������jk3��ݷNp���~�f�<��5%X����a3�6�-�O������_��������I�f'-�a�r�j��a�B�x(Ե�5�~�'�Na��aG�6L<�M�N�O�{b�`VY���@�郟�V|���/�pѥ(�P6ђ����9������`R	T��/��स#��q�Z�B���9����ONp�^�O؈f����@�j�3{��HE-iL"!S�̫l�bס}�V6��3�ڮ��Sm:�VK�0�a.������<nI���M�Ӓ�f����sz.�����'U�y=�$-�� T:�.|0:qwbMN���Î�4��������y�g/X��������)����S> �@�.*p1�Z��C�%}�\I���Ѽ���;u{|e�U�ǶyÞ&u���)����F�m�IQ`�J1G� ����-�=?pK1���❮
K,)Ӂ�Vף	���������VR>�Z��n���mK�C:�g���}*ըz��9�@��̏Ef0��1_��1�j�.V���{�U�Ǫ{'�~V�nt��]���-� 5��ݒcm:s������~V�}3���f�؍�<y����Dy4�B9T|��Ҽ����69qOu:}�c*������G#P�9dRv�z�W�
jLY�$�6�RRR�?-_<�8���<��Ԍ��M)��o�K��l�N0�GtW��[`ќ�7�<*�"Bt�}�_��=��I;h�����Zlnd�@��	��r+*�د5���V_V7,a�>�^u0 ~Ճ�;^���e�]�q���������gϦW`��^�'�J!�Q��Q��UBV���&еD�r�P�����<'=~����cS�n�E�]h����C����B̊I^�P��[n��x�p\�b_�
��kcz|q���`O���X��e��E���E�iRw�U�}
7�5��Eu�é�n���0d�^�g�{G���-4�;!%̈́؞,2V�J���N&iPv�'�扥 �HD'��J�������){��W<��^��f�L����@�m?�1^�9:�~�����I6�;�\ai3o;//�k�,4�	���_֮��q�5���!66H�)�e��}۹�&N�^ڐ��_�u-���"�� #k����tß����,��醡�l�{O��}-�W�\��%�H���qk��À��Ο:���fB�ą����� �v�=3M軎/]/j�G��95r���t?%��{`�/c��&i����Ssc[,�(�k�%��؄�����MD 	���LL�9����q��]���������m3t�_.�[�j.�,B�X�Ł�����N�s��׼�y�)ׂ���E��Q�V�Թ_�=���&�r�fZb��Q:Z�� s��e;� �Ju���RPz�<��=r�ֆ���s�w?����-8�����Z�M�?e�����RdU��-�~ߣ�gs	(��t!��=g!�V��%SY�G3,=|�6X�>{��dSn�D��WNO��8�|g���qO�j��
UK
K\���V��G�q#�F_ �ߞЫ�4�
���{�*]�(�'�Rz�gqW���w��o��-�̉
�$�op��jp�%l�E*ްx�Er�\�=�J��"�����3��=B�F:�ʠ��粺��b��B'Zo��6�Q��{��.��%�	<mLZ��)w�@�_j~�P��W�l�Ѓ:Zq�+���.X�=�)��\�4O�ŋ�C�w/�4��,�y��j�7�M��.��>�x(y�e���o�	y�֛	GL:bt�s-����eM�Ġ�.�*p
�&g�	�h󳙶�{�ܠU�N�����7o��݇�����jOW�1��J�Kx/�����o�Ÿ"T$���Q`�C�`�̘���-j�%�`z��P�y�$�� t3��]ʜa����}�RT�E��2#C�Z���Z���˪s�ථN�:�(�~�,.s^or��o���_A$�z���+�S�N�����|�6Ƹ�� �]�zx/`�
�~����1iU5=�+����\��vbzS�_��a��f��ʠu%�8��ӏ~L��y[����9��z����I����)_��v�:������}�a��!�b��P�Gk�ބ$��ţ����%����
��f����b��w=NVa�2��Ȼ�9��v�ѵ ��ng%�r*��ղf��2k��/Dܷ̬���F��|&�ِa�B�n�}���\��8ƪ}����m3J�K�,�
T�<���Rv�K�e]&hS�_&Y��ś^r4+�{�B���?zХ���7ƅ�Z�B�P�n�f3/�1��b?>���P;h�2QY^�]�4rϱh��7�)�S3�v��<Bew���sm���S4�|�f�Vv	�^Z�ؽ�}�����5�~�_yݺ��la��)�D?�WD���9��l:��Mp����B�%���yA0ى��~�`��дV��A��a?9�C����8�I��҇섩��O�'ߺ\�|A�h	�g�ig�O'n��\��k��U�-�{O����Ll._ֈ$� �����n`�\c��^�`�_	��;K�Z�%�*4�B��+�FH��'�z9Ga7�T�e�J` �:9[��*�^��%<5�S��(���3k>$1{Rl$<˻�[�m���<�{�E��sdU쎱:�T�&5ڭ��c�s���9��;�p'��	�~O����#V�+���h��@qm��K�����8�̻�3�`B�{��%UG!�F�Ėee����^�~ס����N,�H����͒���/�,eLx�%�[蓼謚f��D�^�ƿ)�G��i�dϙ����E�y@��ʅ;XI�V�wj)�jc��ⷊ�����d����s�tuuݡ.my3�b�D��Nm�Z8�Y����}5+��x�;6q��q�|L���(�+Wg����+�/q��p��d�}�鐥�a��p��Q���WT�����*}~�i$f����)�J�8X�DҦ��mu�[�{1x5�$�y'6���{y��V������&�H��I��u[�=r+_����wfn�4��4�&��v��S��H|"��bf�l�b��9c���-��0�����÷T#�>�[�ʯv�6��亁�Hω�S1߽w���]}b����B��8�X&M�JG;2��5���c��������q��h�g�I����>6�j�fէ&\ �A>g%�O�R��>p�ǸV�HY�`����̶'̣��;��0p�#;׊�B���{;�X��f�E:�ٽ_v��ǩ�̃�M��_�yR̀1v��x>ܶ%�J�I �G��I��ۙR���N��.�"؏��h��ef��>Q���$�l.o�\`�3ٟE�|+K�nY@~ǚ��}��=;�����>�$�8H��.����~	'��ej���Xj>��~����x��{�\��;@�^�k���=�7��T����.�p��3M���N|�AR��LT\�54�
s�]�C��e���(+��%4�F���m��:|�(���Ѻ��;����n�����ϒ��4��|%�)������ϼ>�:.�h�㺲�ZͰs��3�j��������{��b��P�Зb�u�Ibo\F��(Ip���󺺄jv,*z"H᯽:�x�&��W���mB�EU�;����ݛ�"�SǦ�7K^��Cm��zw���Nx��Q��03lp��$��G[�1zn^VH�=���[F)�n�`q����qG�9������w_������c�n�v%��N4��Þ���w�3*9[�Gj�G�_���i����ι=�Q��5#��`ăe�}_q���� 7f�/�w<������k�r���>cC3�t�9���9�o��u���bϢ�1V]ahl�3�i3s9��N~�����){=�(⡮���#�~��*�a��F����M�G���Xt�Ø3�|�ǌzG�r�9X�͑��CN�܌�~�R	#�	R�xT�'@j�	������V��Չ���%�H���{ͥDB��8ߔ�1O���_~UZa�&��z���x�x
N��H��%���ܑ'���D(u{�b5�LV�a�����s��B٘E_�*]p.c�Ŗ�y��כr� %���]�<l�o]%�'��6`s����Z��#=��2A��>�e����L���B��@A5Ab?.Ϯ�2ĺ�b�P[�xs+'��R����MoIi�E�ͭ�C�/�'��@��		
��转��{z�P�o��,&l�;��W�s��0��-�3+II�A�L�H�����p+����"Y��]�����˙�q�T��h�.�>�{��F��������"�kk$�L[���$����>(�h4���gI�{ĝ�ȭrjh���ԡ�\
  �d%fbq�*���0VF}g�� q��J��n��I5X�o�&o�QC�A�0e����:����-pv�X4�uN�/l��� !�׃[�V��4G�R�g��r|��܅u���2�����Ȣc~�+`�牀P��_̉���WӞO��%���xe%ά{bV�X"F��&��%�wS�s��Ɔ����{�����pb��!��W�]'��}1�%Ѓ'�&aDBE�'��_�B�d�58�=��W|�M�G���0������x6���FHO����I�pUf�j�6�r��l,�Zq.���o	�X�y}��4��Xe5
i(A�A.f���$�Wbزm�[�J�ʤB��K��=��xȃ��w��;%!8]��qT������❯f��.�g}\��7�b��)w�4�^�}ї�>lh�
��R	V&�T �w�'gm&�4��Er�]�����ڻ��r�dh�f��D��a�y��uJ(<��z�Ո맶ȋM%#F�����xĨ܊��i����t��UB�� A����9�#���9���l	>��{h�����>��r�a���v���	g��� gg�{�/NS!oǇ�*��qY�$,݇,Hg!��U6)�kJD�na
%!W��C\wH>��ca�?��Nǂ���kz��� Ph9F��S^������c2�<y���(�-zm��q�6+O��Z�y{
]��G�j
�jD��'�ά�5~-�J'2�%2;�SQL��y*�.#��p��)qH��� ��bK�B޼g�\k�a@i .b�,�0�Nt�(�s��Dj� b(L��T�ʖ��y50����t��}#"��]�������1Vi?���4���D|rn�-��X�]FԊpE�x'ki3ڀ�fh�C�����(�W�埣��x۳�w�Ӄ:_��bC��sÁ����oRY��	)�4N�t��X-r�>ن���fP4[����E�Q����H}�7�&Xު�)��!�:k��,��KC�,�Hu	/����򀀌&� ��a�M��SY|m��y�ƮT����w�� �}J^�R�����Y����1�fΔI��K����M��œ}��d�.����ӫ��@,��Q֗�_C���b��w�a�o#siJ�i͂���S��'6h�ⱳ g7)���p�&/ ���`s
��<܎0w��c�p0h�h�5Qi_/̸�.N�v>��l��M�Y�1	�Q��u�/U�*���� �7ak�!x��E�wB\Ȅ���$TB�-?�8c�z=����ZD���B���A�+
~�Ϋ���`���
)�3'p�:�k����N��bݗ��u��}����KN:'Q� [��I��k۴�
�u������E|)Z��y+������"���W�q���6jl�7��=s�^H�ڠ#�r�T����B�{���:���H�z6tn���ED<dB�X����}ܹ���y���ku�bSP��.rE��_Z^5�G�x�̰��W	2����6i^!	�)[�(/�Ѹ���� t�t7�'�>��zIX��y5�[�uW��"��Wn��屁cw�C7�Q�7�%�~�������������� nA��g'�0�1�h�mS��3۷���.�A�N2l�՚�Fl��@f͎�W����8�u׺��q�f@��%�:���x\���d*}�o"�������SL���u��:9�­��:NL*C���ڮ;/������������[����B^����a�5�R	�.?���o|��^��b�$���h�m`a�*��H����PpX���ۦ�g���/�m���b<h(���B(�؆2x�輹^s<��u�'���ow)Tc2���;� ���I�y����K$��yEz��(�qY�5�11�oH�:�M��j�B��7�:�^��k+�g#ˇ)��,�b�Ȋ]��v�,~T�3��<��~��r�w���F\;��﫟�ܝ�1���!̫�S�J '���N��NO@��mZ�q��%r<�Oq(�&���fki<qdV�3�$C�V���5Ig���Y���Zu[�	ў���®rZ�wm���^�xe�����U�Ó�7��ԁn�)k�ѱ^؊y�vm�^1��)V\X��Es����)x�
RNcu7*��u����ő�'43I��b�ם2�}F��2W�y��@<�ic����>N��f�2Y]��Cz>B9��jP���bW�8��- H�D�
V��VS��G�[���~��s�/�����&�^��[�鈘���2��=�� Y_q��DY�Y���G6��Y���QM��9�(����'��9�xf/U� u�.�Rdk��m��k�R��,D&(���]�� H�[��s�
���O�__ �o����
�jxQ.��n�\��]z�s�@5�]t��ۉ����=�B�{���g5+:�<+�[�g�Z/���o�t�T��O�	S��Sǆ������j~K��G�W&[�.��q��#�^�ǩ|��OA�5�� �[G7�&�t�#�yW���Q"�/��{�0�龖���JS|d@F����4a%��|������zzA|q*D5wat{}~��?OωjA���-2h��6�� #�ɖ�׿��s�H��_�ϗ�g�B���/H�F�>'�I���$�i�@���7f�@��jED�~���"��1�qLX� ��R����~��<�7Wb�+� ٬u*��FLC)�?����r�� ���	E��x9��>�;f���a�\m?�$�a)����V�|�Ġ�C�/!��pC����X�B ��E�"��JQ>F��f3 ��cu�p%+~�2|p7`�J�ߜ��~a~�l��;�R�ul���6���	�{�D��[���|��-�Ue�rBAB�A����0خ�K1s��4$ ����@{�?= ��NŃ��~�'߃`���qa#X/tTJ��1aP*�JA�+b�m� B�	Tʪ��>O�[��_��S�<�b�Z������c�m��::���B�}`�ً�.1Pc�V��jd�b���$��|E� 1ټ]��J4ɺ�<4]�ܺ�	@
���@d�7�t�v�����^?O��tR�����ܔ��t����� 9Sxk*[h�����@6�ȣ%k�F���t���O����f�C#H��kSx6�����ܦ\�D�O�Ɲ�a��[�K^�D ��1$8��N��9�GZ�O��)��X�Y<b�V�ύz5�:�gb.j4�h�`�����`�d��"e�ɣX�7?�Y�D$A�CC�viN�2�n{B8�l����f��4���E*	h=���qQ�Z.�� �!'�w�/���F����~�Np���m�������"��w�_����╳*��*v�|=o_�=F#����0�a
8�4����i�K�é�1e^�4`�KxLj�so��K��J�ߖ��.���JǨ`�

��^fA�������7���-`�$� k�/�'�)�P� �bG��,��v-K��ϵ=ۄ(
o`�1q�GH�]����Gݔ�7�i˛\��
�
���GvE�s!jB����֤�v��ω�&�CL1�QH�F�_,d��e�΢�B���L�Kn�~ɐ��n�%��ZO	�9�)��]�S��r�J�n,E�J�@!�EI��	�h��K&�ԈY[^j7�ݛ��!��,s�4Qt3M�U*��:	�>dt��_��&����$-����셼2ߙK6i��6qk�h����\��_2n�Z3�<��+����'�Gh�����q���m�5)ȸv%y��$�Y�/-*�>��r;���N�K��zc�:�@Ǌg��&��ّ?ު�����7�f�*�fjܳ����y�璡�􏑙)!��h��l�AD2���k�w�&����1�/�P��aCd�� �@���<aG��	��?�9��B��>�ܢ�Ã[��a�9(�,���:P��9@��	��p�|�z͊76�҈$PD��>�B\�2:�w�ȵ��K���G�۞�!���_i5wRYԣ�m ŭ����o�B_l�5]�Ԑ� �&��m��3=�!VZ�cE�����ѓ�b�B�Y���${]#�w���"�e����F
K���JVPƺݴ2�an�J���1|ac
��0Y�H�H�����d�qx[%T5G�� sX[��[�*�(�hi��k[�;D�as��m�
M�j����?'��a"(�@�mTҘQ<�.��<;f4�g'?B������	'X	��!��Q� �4&�)(�O����٘c���!��*eJ�%��dkt#Y4}6�H+-qҺ��f��Ǟ~K4Uq0:���=�GrZ&C\Ȯ���K����u8	Zˮ���m�I�IU0$�N�^>\��aYrd��"6F���[�����9����ԛD{˟н�KcX���~�D��78{;�3�Q�&3_��0�w��cS�Q�Ĩ$^H�!�s0��%<�K����
�j.5���c�'����+��~����g�W*��o��,Eyq�@B����/�_I�Ӫ�i�g��c�����?l#ϐ&͈��뜕5fN���M�\�t;��z�E�ZrQ$�� *�؁�e��(�#�l�,Y��z��=^��4y�����3д�%�ޏE���8�"�I%6��}VQ�9�'_xh�� yD�Լ��O������d%<�:��Ơ�~��ď""u��X���*������>�DYW�GN�$
f����	�ec���;.v'��㺽����D��Р�A/t�W��&�M�#@�"R4FN����2�0�ra�p�j���Ѳ�I��0ʺ> k�;[ք��+0r�FT%(�v�-���;�q�AQ�� �!+�8*�"�6yj��:1&�K�,Bpq���J�FBM�o���δo���@p�1��i���<���DSB|L��8LR"�ABw��~]�J�vh��r�,�խ'���G�QQ��Y�%P�
����k��1��Z��"Q	�Nz>�.q���3FJ
ja2���B�(ѣ�=�$��s�0`di��pm���2��+����Y����2s�J˓vmH����U�aRR0L�Ӑ�Z;<}*�����^�ƍ�1�Uо��J�c�2H����F�Qc�|��} *~�P	%��Kt"5�+��I?�(�SP�0|�]q�>2j���&�|�!.w�� T
��B׷ �Ȅ	�S����"1�9����,3��{��>��	� �S��Mi�1�� L���7��5)P[M���9Gy�a{�B��¬Jh��Sy~�8+�͉-����>�@�!a�7#��[�0w�(��O%+�h<�)ƹ��ɠ2�mO�����v�(#��ݘ�?0m�+��|2c�dpt�y)�&�!H,�s �7@�hbz�¤��t�BF/Ch��F��po�����K�.o͎��I�_��p�BE4Nq���q������A9m?���H3����l��?%r��o�*J+N�*J�{�O�8��R�Z6�"	��͢�$G����d���+�kg�
\�
L�n���Fx`xt��+��ݯ�~��u�N>�.3hm�)�CY�M>O�]^�> ��r�)@�;,͗X�2ǡ*�Ƴ˸����rf
�&襳ן�����%+�˞�:k� �4�y����Z;�b�Ve�����sT���Ul��D�<E֑��M��1�_[[{\.��Y�'v�$
a,h�5#��5!�{q�dn�{c:�]V���i�|3�(AE�R9X6��ƀ��"Θ��6 -W�D�����%Խ�ݭ
�W��ȡD�"���KA����[�K����U#�/Ն��+��^��re���#d���ö�m��2����4�_6��_���
��Yp�{���	<��������Q�p3��������qF���9� ��k�:���y%�J��#`�:( l�'p��R��P���<��^�M��UK-t8d��C�����_DO�6�5-2!k�����p��0)5R�y�M|�hCu/Z��R��0*Gv���H�ly	C�3z�b��A	o�<�a� G�:�u�b��]��P`^��񋅚��%5G�9��?,� ��tD���mb|QvN�&J�p���:�5��I]Y:`�8�;�O��w_.�p/o�h;�:x�*s�U�^G�l�p���I<dd�?+���Z�x�mG}���;\۹����v�X>�׾/�k����@0��6F�m��g�/��u�mϼ����Ȳٲd�{�R��;�Y�@�M�$[�~� )
�<:,�d�d�<����^̀T�$�"��{�,D�,<�ijv���(cRm��3Ε5�H�fƔ�L��O8'����Z���S��rc�E�ͷ]��H5ܴj����F�mMހ+�Q���23�5�������'ohʆ�RP�6(�E	gB��B���M�s 4qH�T�`�D0`L�>	�
��IG B~���Qc�!@�v7 �
����!vb���_X��:M��w�����Z�4c��/QM�Wj =��ư�jA9U_f�@9Cy���I+���P`����|hc>(I$��Yoo�΀�l�x���I4� �싸a'~ȝ��'C$)<�Vѓ��%3W)^�i��b:�O��_i6���)���}p�Ņ|R���
oX��-���ޚgH��� ��pE�J��D�Y�@p�ƕ)�Q�XENl�h����rH�`k�5bR��9-E� Ր C2�8������/X�C��]L�
�PqF餝���k9ׁ{{��>Xα?{�׼��N��$>��� �Uz�+㯞b��Z���#+��]c�ˆ[�2��y��?;]����=4��ǯ���lIcS���?u�y���{��)x��S9F��ո�	���,9�^���`M�
 4_G�DLݴb�Ǌ�>�B�ۄ-GfyۇZQX�!J�B�Br��~�$�TF'�e��<\�p�T�7�<��%�y����0��J�tz�$��
�+?S/*x�f��ş�%�b�8CZz��;\:/7�Ql���]�X��l<��0��;q1��@X���f��Ƅy���X�f��1�'k���yXBm�6Qi+����#�Z�
���T������\Ï�~�8�*Ĉ�<���K�s���.̟vI��l���2=D���
Ka���V/�4�*/C�SgoT����7Q�C�]�;�ø��l�o�~*Xf�	�G�/���=�:��7��R�o��a�Q:��mc�x��f�'֪ż�����3H��Cu0��l�J��~9��A0�M���t�$z3�gG�P�(�� �ܻ�^��`:G���nژ7+k4���L��	�b{KT�j�F�� ,������ߥ	˫u%��Cy����:��Ǎ��'�c���c9eS.���	�?D����@�8X)(��R�,Ov��N���f�<0��
e�������F"�z{��Yp�>�F�H�������:b��5^�u�S����1.��!ڢ��G!a�9�B���N��A���j��&s��p�kM��X%x2K�ӯb*��W]P�c���d�� 3+��ε���u��8`��ວx[����b`�!DHQ�,=(����j+�6��������/o4���btF[�6�dm��
?9B >i#��;����|�psם�<~��Y�t��C�A�=B�o��/	j^�I��j�yN@�
zr�$U]���{�a���Rm���h�6���^�wϥ#�]�ؾ���@{=�=:$AA�q�'���(s��W�u�%8ǽD�1{��_�fl��9I��҈"�M�����jъ��6�p���{ n�[��h1"�z��$���67q�AU2\=m��(��,\q�����r�e���ܸ`]�-i+	�9u5$p�^'��9Ӣ�������ӡm��F�6t����v-���o�_�惇�����\�u@������m�D����W[�"�yد���{B��$�������mO%��l7�VW����BG"E�ΨCv{�h`Q���4_��wx����w����]�0�Ed�����M�oS[�%.j,�\.V=�8tz޷��k���*/����m3 8!��a` �xrN%n>�������R2�d"=�L}:ZGV� ��I�+����|�1S���O� �O��5N�|���r+tnFM�U}�:oPR�3Ћi���R���z!^������NWomh�����"D��(ԌKx����Gg�'đ����t�dH�F ��=�������״uk���J}��u6��Gb	ĕ�5���!�j�c���}��䶽[���fΞܭ��S���wG7O�(Θ�^4��m���	W	�ɭB��Cf�	�F���*j��";��ѻ
�������+y���sHF�kśH��xF(�Xh7b�^V?���-c��<Ʋ�9n�9��I��@���YO�1v/<��hQw����)��А�}���;|4>ɜA�������!'C-�9ݺh�7�O��j[�R�Mer�r{T���Φ@�M��Pi� A"'j��֝�f��F��k��I�;0HH-���%���O��*�04G����Ī:C���,E�34����y�.�0���ݦj�N����e8�3ނ��_i�UZ��V����7����A����2+p$)�H��v�S�����{�̸�[�U^w���^��yN�"e�m�áM�밦T�	� ������J��������pf�p|:�W9>�-�6��4n`�L �ޭ�$����'�1�L�)�8�un0Xނ�2Icⅱ���xLA���YA�zش���`�Ҹ-���߲���u�CV��SYcJ�����/h[�v|�n�4�1i2J��*��"/]�y�'<�qQb���ٵ�ZT�@M��G���&�}΍<7�sW���5M����']��{�>�U�E����n[�^j-��t��o�v�ww蔕X�\��_h�]�L�vⲾ�t�;�~,C|��b��=�qb��h̾�2&%�HD��9Lgc7A��Ch2�f�c?ݪ����dԸ�}�Fʄ��*A}��wIO�c��-Ěf�8�o�3I)��ʎ�(]��?o�5��+�~K[�Cx ���!n�h#^=Gu�����>s�n��I晃7`�!�]�$�{� Q��{���s�����t]=��A�P��?wZ�v:p��^نn,�����'���=����f��e��_/���#�F����^�C{!��6�6�۸%�^<n�l��aTv8��F!����}x�hva,��ЦZv�0�����ZK�*V���{&q��=k�b�?z<�����Yo��E�.��n�5��C �wwwwwwww��	�Npw�[~���{U�j�jwg����{�=�g��?�M��(0yK�1�Lv��*u��E6h��MuT�7�*Ȯ�|ȕ�Dl\�G���.w2���-S�q� ~Z����|Lgs��n�ŷ�:k/��G�{�6�	m݃�Kqs��K��I����$�O�l!�B#-��ă�j�y�bP_�a��.��K,��d/l�2��6�9�Qa�㉜��U���/h����l@�%�=*ZK��1W��V�ċ��2�����xE|5��<���)�-�\���=1��}���M�9���k�c���E)�7�V�U����N�9��Ӻ�_�l}H14�5�7�MU�=�8m� -�T�\�J�R�-tA�^�\-��%��..�/i$k�7[-��<�Q�
=�2G�8�����+�>�?�{|��(_l��xU�辆LR���W�����T���@�׏�X��0^��lg.x�����o[jp%uH��!��x$�S��1z�p>��ce�ٌ�k�`�B[r�8��Ka�6kFuD�����.��
e�*E˟TK�#l�D�[����R��Ƒr.� ��Qbv��*Q��P~@��>�d#��yj�~a!7���&�wܵ"�q�m�ڮ:Hg������N���m��'l��V���G#��%dR�呈�㠟�b8��`�̠�Z������Έ�9q�ݎeJX�Q�&�u����au�#t �>�P�ݫ�G�����ި�Hu�N��܄�]<�X�ӄ#�d�ڋ�����o�yL1�S�@Q`r=�3;,rH8!�� 8�,�ُ5�٬��}S���4�,u��^�]A%��<�x�캺N��x_���V����~S3�=X4�`�j{����'sm����m_1��H�UB��Բ]v)Q"��6���3rLr_��p[��p��������BK!�&�K�����wخ�Ko�ٜ���FW��(���"�b�s5�-֢�S��pc����r�r.���ɯzX�2���#��j��d���M#���"H�#��U�Fh�H�ZkJ�_��ߐ��c?�Q�;M��=�y����>"D>�y�� Q:J&�F�y`o uf�L������~>�~��Q 0����͎�_�+����bP�C6JI����T�q���n����u��q�m��j/�?��l5��	��H���a�z�)�q�Rf���iR/j1b�#��/�ׯ����C!��f}��4'��亵;���^d�/��%�X),8,����Z{f��IL���)�����Y���.r��[o�����>'1'&�0y�>���ꕍS<,���?�B�VyJXIe����U�`%69K���t���b�PluUsD�����	1!:���I��� ����_s�;m�3q���X��,"T_�.->`��^�v'���.��Vq������y@��y�0B�e%�A���X45&����iV~�g^R��WZ���t8),��$Ðӷ0ҽo~D�6"�����O�-q7LƓl�;��?f�c�ٝ�[]��[U%�W%y��U�� ��<{�V�ǣ�/J�!���.���|#����kp�rON�}��"3U�#�Ms���|�G�r%��\���	���Y����^P�G�%���y�|Ք/v_:��im���{�iV4].vZ˒_���yc�
�D�Zz3e�`�vY"�bʣ��9JB�E�<�H^�F��k����F��)�@E��]jf��(�+��58�'��'g�R��������Wヂ��?Fz.X-C���N�O�f�h�X��H��DS�y>��hbv?��8��2���g�i�o���)ے{�B5���ds�8 ���)�8b�\�U��|��a�J��7#\�I���C�1.@ߗi�M�뾬A�Y�׉�$�d˟�zܪ�Hߦ
EJ�rIa��J���b䎦�J��a �F��Z�ʪ�-�)d��5�(�W��JQ�P�͆���uC"���G!���{��E�f ��� v���X����і��8vU�m�u�Ʉ�󴡜�)���ΰ�Fm{BC��ܿ�e�?��%bSa���;��;r�ГqU8�� �2Վq$i%��qj0�<�@-5!��}��!�H��U,ۛ#�A�/ʛ�n1=.*����]��.�R�ٕ��H�v�@��b���#��� �����'v �%PCLk":O.�_�7!M�p
�(�h�s*��eH����p��Xi���D� �(�h��E������[R��=c���%�oPzb���b�9�K��L�d�-=�^����b��@E���T�ͨ������K������24�M��
-ǝ�,����o�B�.y�Kvv��8F!I���;�1���{��q�.�+��z��oBZg~���*\�ď��V�76�X3���#�צ�[���Y)+��"�Y�(̎����_�Q�u.��Q�b�:59�jM:f���#����0�����J_*
�xK� �$�`Ie�Qq����yV���f�"�#�0�b�#X���_���n���y�k�O��	�v]�V-��j�S�rf3`��R�ԚY �耱��BN\FR�D@ӎV��]V������ËVR�+�Wa#�Z�W�����v�
�g�3�Mi��%e�'� ��Pm��M���ۥ��������F�I_pI��~�evX�4x���I�ƾ��oK<�F8��Ҵ���������~�feb�
�0�s�I�Q"�}�x����e��T�'�wZ���~,����u��l}oh�>v��������2�bñ�G��{�acMu����ULw*z%l��bsd��� s4��7���ƥ�q�ُ�&�[{���^%-����������^��s�n/���.�$��b��%lG�?)sOh�*4�M|�N��#�KXJ\�8X�0��5��Ѕ=�{�]���"��nfJ4��� ��L�(��#D��9Hug���@(���jׯ녔�#q��v��HhM9n`i�����n����Oi�n�w��'ʛa�}3n��N" M(��3��6�L� =�P��9���n��n{�?�7�Ȓ�e�C���c���i���E:b���)�[�m[qVE�����cjd7�G4��?g�v����u��g�E�ƔV�A���>0���oT�=�_��|bc��@���&�ѹÍ)"N������7S�n:�;��M�ͯ�mndpWt�h���]f]�����
2�?W�^g��øT1V��τj��;��Hn
��Z�P�&��ݦ3�p�8��t2�5��M�haޅu�Rj��5Hy���.��^������h/��Q<�<��\�ԓ�D~�La�N�F�� �������vmK%����-mȞ�ŷ����8��^��GN�2ρO�2wV�O�4�qFH!]^�
@�83�@)�G8��8�K�9�̦��s�ӓc,�_h
Y&���P�=L���um�ZQ�lo79��|I�||!�QZ�T�9�,4�5јVl|��T�y&I=��|1k�%�ل0S�"c��~�+Ľ����|]@��+�N�ã�~�ӄh'����	{/�.���|tĎ<zJ��J�m^�R=���e�Q���z�fg�Bգ�:l���X@-��JP�t.�*>�8�����}��K�D�0�,m_��"����l ���9?|�'�9)�%.R?���˙�W0�P2 cb�%�dm0b��9�l���O��@�,L��%4Ɏ���J����\7�E�=(`v���lP��Wu�2�S�Y�Ğ�lֵ�8���:x�z������*��S<� ڱ��agb���Jv8��s��4��Q���6?"d].���F�����С�|�[�)��H ����r�����2D�>�FѰ���KU^��I��h_QRE�9oO��8:o�*l��ͭ�-.�w���9c@����RL,��.d��$h��J�X�na8�1�Z�9v0�^ى�?�T�;F[jc�l�i0q	��(4�3����ߣӸ}�J�y1>���W��.�����	�#^�����똉J5����&�4`���~�e<@[5PE:�	�^ǫ�~ŕ�c�?E���p'T����_Z�t�@��5(e�٬��JW�1pg���%�G�}h�-U�X���af��q�b���<�-���[�=$�
�,�����+��+�a��q��ޏ�g�;	�;&��d�_p�4tx���F���2ܘ]ʫL����}�wN�<Ԋ�]t6[y��Ȑ��9R>`�����7��H�d-����T6TǀҾ`�&�����|UKsy�7}�I�7����Y|5�{��9a�x�p���*ineu���׶1������#jT�������*~7~j���t>I���� Q��j���7��ō9J�u>"D
͇����0��� W����[*��߈B�+ ΢�hDx|��h�b/ڑH:�� �nCC( ]���8_A:sGH���q���X���l�Xo�����n�&�m��iL��ٺ1��'-"`.,�c!���D�w�����J�����D��ZE���(��N�*��Ǡ�,)GE��}��{/@�/x�\u��,-b�0�G��_�+�%��]�\7��a,<��e\�-�n����խ���o@�����J�滋H�"�	JD�M2��s��Jx��t�а�]�����$a����-֚R2ʲ��Ώm��i���-p�Y����O��24k���T)�5�U��L�^��-����E[/�W�&��T~�xI]�p7)Y�GBѲ(�o��)�I���^;U�[<��7���P�V?�Ŋ��%�i&�թ���Q��L[��d'���؜|�3�&�=�*�XMp�?;J�Mz�x�m�2��(cuz�جG#�@��f�R�\�%�қ+���-!��[��0�֎�y=y�j�=����>�;y|�v+���-v��{i9���j(�v9Trs�->v���V��q$�\���l�s1����IǇv��0s+�ϮW��S��R^�(Ix��L��m~㟹�%Ć�q�GH'�|0�6O�.��>�e%w
f2�*��K�X*��̮D,Q}��~V�5�����'��2TR���v!J��w�������7:�'=!e^�>^!}|�{�9W����JMa?nJS���P���1�l�s����wKo��UZG�G�=����\[l.-�7��M�q�e�xjj�o� �CiV҄<7�����ќ�K�,Z4K��K�ݶ���ވ�:Z�oNbS�^��#��-[q"�N<i�!b�UQ$���\c�۟�Cs�W!x(��G��U�)a2v��5�cԊ�c�6�I� O9�\�]�QEk��2'.�|��u��wP6a$ƅ8�EH�|^�f���_�g'���ie-��FTWĶ�_��Q��Ir;#�;1�~{A�6)H��%���/�bb9Iϙc�W��1_m*W0��a�&��t��S����Ҭ.C�6��)��oQ��+`�CDp�Np�c��̘�3�tI�gO\}�����q�{��l�]V����%sb��t04�X,
�&�,��ف�/&�i��e �f\�1"sЖ�Z��*l��-[��[�a���E���:�] gr'P��7":VD����?'��;c7<?�k��H�z����iP�J�(u+w.�5�w�6|���@��S_]���	�~�^�o���Ϛv#�kxk������%��A���ҳ�X�ɉ�kK�uGE0�U��~ǧIߚk�tU경����hh�l�a���B��sM�s�rp�e����� ����	D6�;|�yt�l�X��9�ǃ�dT��H1
Tk���F��m��	#{b�#�E9L�a���'����D�:��S,9קϱv�$K�|�V�q !�J�sN��S��%aD)!� B$-�|c�f�'��"x����d�y�\���#Y�����&{�*ӓi���wֆ��\��p	1,��Ѩ~��*n���ЛX�i��[��<ZD��g��iU�-��V�n�Z((Q�A�I�ۦ)i��Sk�N u�F�L�1���
��Tl��i{�|������Y!�;�7)��ӱҳ��4�S�(�+M�Nm-��*��_!�r�z�B�[y�C�2�\��{�#nM�qIv�1	��c����V��b�W�h�&�H-O⤯�3�N����d�PA����+��g���'</������B�P$-�̼�`�[B�0f~O�z�X��;=vKs���k��&�������A֕��*߻�;3�࿺?B�q:���i3��;)@�S�(��쀌�I%҉CE-W/U�����9L�=�'��pY-�����X�uQ$ѩU���E/�DQq�fW�M�m>b���)Jmgs?@��A-�o��
���l�j*�*]>�$eǂlu�ٵ��5�Z�e�n� �"����+{9F!��1g�{�F��
U��`��)�'��%M��#\�sk`�SĮ��}3���1{��&�^�`'y�J^MY��?
$G
�$�'�"b���ha��o�}=W���`�/޸�ӟ<Ae���me�����x$��h	h}m�\�z�;���u�nBCs��9�ޜ�6nU��)8U?�,f݋%���I����Q�8�y$�"i`�^ұ0��뚧^������Wpc�l��5#�&�6B���fղps���qpi�Y��pv���um	�MRF�*P��#�,!��L��GD �	�2�X��e��������o��"�_��J.��Ԓ�d9�I����B!4��qw;����o��ar��($�ĥ���LG��f��UJ�L��E���f�c��,���YrtZڮ_����F��^���B�)pw^�w��}G,:��PC�����m�P�rY�_:�%��*�Tz��e���R1
�R&�c&#�&
Pj7J|�=�,�ӛ����Xy��)3Hb�7d-߽JĹ:�ut��D���4��~��w3��[浻���3�$��bY�ܟ���H*�y���cdKS0~c��@v3��Z��d0p@`g�p�c�#qDSB;����Jk���K������ލĪIO��+�[��M�����E�=5]L�qO�f����v&���,��\&�����&^��"wk_�6/�����'��ݕWh����F�9ոq��qL�+���ܨy�ti���]�ᢐ�ow�2Q�}���t�襏�T�,��ދ"rz���g��{���B�΃�+C�5�,y���k0@0$.
��b�;�laS�M��//�|S]��&V���-�\	�
Ib��Q���"�wg|��x�z���H�w�Υ��;��KiN����������	��-���?���\,�č"j{sS-͝{���һc��q�� �)f��']��-g����(�O ��S/�f$»S,g	������FN���j���u���9W�7� �=hHͤǯ���m�� p�}���`B��W�'����b�t�_>�_�D!�Q����4��νkzI-�L��#�Z~�;)���q�
=��P���%N~R�3J�MU��٦��`q����j�<`
�M&�ȃD���Sk����"q���f���i��tv���s�(0ahG�,����1/�[�����:R�"�-�ʢזk/M�k�߸�ܭ�G�M���+O�3���$�zЕ�{a0�+9E�ύ%B>�~���..�B�%`/:A���M��+O��[5~�[�3��_�����BvOe��e��K"�"m��D⿳甏����5j��g�yƆbu{�����Z�X�=�X$}\�.�SQ-�����/7E���豨5�Y�%g`<�~�y��y��_"�k�P�<�@�p{<�'�m��(�����T��m؈!*6��1�s��U�Gߑ�{�������W�	�qDTf�,�eu�@�f�������R\�{<l�1�<�W}FN@N���D;x��b
���vޘ@#�֞G�s��p%��B�׏�uW7��B�����*�ƭ��KC�zeGТ�Ұ���۩�\�A�E&�)_2C0dKj�3��<��*Mʛ�2ul����gJ&��b���o��֩��:�.x��!rq��:?�+��ä��\̔��ܯvɒN]��Lǝ����9Y  Z1Ls*2�m�)�J�{7�|����~����f#��A}�������nh葅*:<�Q<�g����3��j�v�0�ߞ���_-o������t1��P5fW�Q#08�y�ں�����'�����b%|�dz���-]���A��ҳSgɪ���x��G����]�=��>#�n������z�Y�$�$f2jYؼdTk�j�Ȩۺ�>��H��Y�z}�'cv��S���Cbr�0c]��zb�c�S{}�Jq��R���8s~'�rg���z�_B�_&eϚ(�&����k�Z(�'�L���e�yND��r#sf"!���.9´�#������N�l�W��0�>j*Z̙��l���|$c��.��<	#�K�t�%�]�w�W��d6\���E�!h��cQ���+TǱ��J��)g*�AO#߫)@�F����#j��Dv��8�1�#�������
���������q ���C���{� �Ĝ���mT��N)�bN� � u��T$h�TA��!�O0�>;
m�l=�+9o��i	$ĺ���L�9X��]C���!#��U�Ow`���_��u�1I<B�G'h����j��ȇ����������;�y�/�c��M4����D���Wr-g���TOT��x�Wqɑ��	{O(A��a3�\�to���F�l�d�)`�/���9$�1Sy � mؾ4iYzѼ� 2�N-U ��v
�� ���O���w�G��O:,\��z�|���������=�U��W�K�?^�N�9��&���
̹��D%�.ѐ����-���r/��8��0R�e�����3�t=}98)�PY]tb�1��K�U���&�-F��:YAyg&���'�?_Y�[�C2-;:$K�J)~`�SN��8n���Mi	���%	cA�����
�y���?W�B�e>Uf�t�({�����d_�\ŬI+#+1;��fD6��Y�Vj#��Y�L,Cf��/YCoȃ��P�5�AJď���<a�X�����Ȭ���SN�L��z�1r��&�p�3d.dm�;�e�_z)���?���<�S�嗕�b�/^��A�geM�R$D����1�Ox�!��3�#pKv����aT&;��U�c)޿��8/�����%%�h��|�j�i"��@#����槟�ŭ�
	ꏜ�^{BHaRԸ��r�ɼ�{qq��hF��/r>��~���.��G��f�G���L�LYk1�qY��g�J�LS��u��P�!pL��_{�Ĺ�P�ٵx����nL�n#�z?��q�[/�Z���*�����"�c�����e�]�{�2�ȂPəE0����,5/ϲa��җڌ8U�L��6��W�2eM����pG�3#�5�|X��+���"O#DôZ��5��pk�(�0�e�����0��M&(j�J��䪟�k?�����dْ�ēz����~QT�͇�������P�]R)�;�P.�nν�ϻ.��Τ�{���0v���B����¦�m�a;#��T��=���͗�&+���ݷ���w�8Ʋ�<<מ��41+��+{)��z*~��ASJ2䍄KV���JJ��&m*�9�ЂT
8  U��ͩAEh|�e�Pj>����OW��9�T�}@�\��9,�t40ș�}g~�p�K��*hV�)�$)���>>��DC���E�@�x�gE��1�X��s���i�E��ؔ�6˻�Iv�l&��r�����& ���筇j�k5�Ъ':����-��o�P�g�����c���e:/;Cr<�#'����w�=��H��0�L�hJ�~ ~���Qo�)�Ջ؁����?oMtDx�1���g..�;G�z1�R*>x;�u}�>����歐"ah��[��x%@a����|�������(Ll ���/���1izI�!�4�:(���v0�h�����ï;wU��{�6|���{�Qq׫X�q��Z�m3M��1k������P[p>�����V'hP��(p5��Q���,�� %��+����&eg^��������L�Gw���X\
��)�q��r�O�$Vo�������'�4�7˂e_�ּ�_��2k��-�1"D\�)���
��X���aq+m�(��u+]���G1�*g[�k5W��^�������;X�ͭ\	I�@"d#Z��4��K3��
��Q���U./��Iw�e|z�eSl;\������x�:K���J~Td��>���r�uPuh��ד�_1�#�ƨ����kbJ���p���" ��t�PW���u*�&�I��4���E~z?'Kǉ+_>�߭x�P)R$b<� I�
Il�´]�������p�:�[���������PM9*a;����z�PRD��>�਀����=���p\��v���N^
LxLx,5�����G ?=?1��$SK� �ګ]��*F�l����ϊ����ˡ���]���������~9o!X���Je���-��M40ޑ��D~  �VLPL؊���WH��i�F��hX�O�=�K/ �A�%��Ȫz6^�R��q`0�bd��ۥ��x��b� ��Q���<�ta�N�qX���H<�E�-�t��L������F�J�}�<�0���%�v�8��v<ѩ�"��eZ���@C.O�������`6d�[�� ( .�����F��%��'ؒ����Y��cs�m#EH�/�^G��kik���ʡV�1HmZ2����k�����^9��x1�"�˺�~���V�Um��ڢfG�
�A��(�D�__B]�U��u� X/��������nb̌��H�T�P4�+Ѽɔ
�e����fz�-C�K��WSx�qh�儚��m��0�\#c�&:cZav���ƑL�eX��R�_8�Zk(�(�MŪ��6�#�q-��~�����	��Z���c�MA�y�E3����E�V,[��(s_Sf�ik�2�>��SA����cg���E���ݍIU4������e���\� ��_�Ѡ3��������%S��T<�(A��e�����rG����J����i��[f�v�0:�D�kE2���m�F�B�m�K� K����B�x��x��@�7�g���ŀh �2��πx�`9b�	3$3#!A�xi���Q�f�'�@r%����u�#Z�cƔSH�n�"����#{��O��CVB)=`d��H�U
���d�����&i�����W��F�Hhp���)}�+���B����9J�������Y�>z$�;���IH�(��tc���^ϊ(��k�A�[5��:�b��)������ ��mPI�g!����i�	� Ɓﭡuud7X����Q�Q6l���� &P0D��k�1Q�1�ݠ��#U���/��	W�4�~���|����������#0��]I}���~22�8ZN2��2#q��|�P9	��=
�H/����C]s���O��WD�;��B��f#�ϻy�ʳ�r?\�ӻx�y���&���pX�#���ٮl/�cW�O�?xF�֎�֮l�+I�+ǁ5l�~C��|׆�zX�jF�CՅ���?r�?��$�%��[%�ȋ@�zbB^�L�����(�$��͛ޢݪw�@�:߅��Txa�p�����p�a�XwJ�R�':��!����Sb����P�|h/n�?)�5Cd�,��Mb�ߠ}fŊ,�W���H�|+�0�^�:�;G������Waq�~�_��/4)��E���Ç�Aq��5+Uho33��$lt����S��|qFJ������9����[O�g
T}��8h��Q9�P�/Q!�Z�י,ĥ�߆��A���q��9��cbs��#U�h"���D�5�����季47i�Pf��ry�L��-���y��u�gcN ��R-��<2�����-+�K.
�������m�p48(��bwkw��/E
�b�+�p�tL����,uP�@�G}�LfE�"(ѽ��9dm�7;�s=�bD?�nD��f���6�L~j��n���{�׫᧸�.�uю�`�xΨ���`oE[$�����v�ؓ���r��^�ʙ����<ݩ�1X�ʐۇ�ё1��a��M�r�)��=�7���eOj�_�n�[qVcR���k�"�'RS͆^t�q���6������F5��Ϯ���z�X���f��l���e�f�:�>|<�?��{�|��k
 ]#�a9��F����GBKb+��h��L9��x��K�Cػ�������2�<8Ć��y��u�^�~�7���5q�@w�G�d����;o���oy�K.��1�}X��QTh��Jܲ���j�H�M���7���-$|��\>O]��(���ܽ�7�2;����y�<>(m�w��l�� &��X��V�$�"i�c��	��K�Pt8��5��5���"!s���Aqpb`�}r��;@���Y@����T�P��ϡ�j`[C�_R~�4aG܃���n$�/��������/U����W�߆=%�-�B>O]�����<ޠ0�[�.X$z�`���>�XXx�Do���0����sx��T����zO��f!�/�VoC�QZ'>��5�;��p�����٠3*L���Y�Oɛ�/h=�(b�GHl"0�,x�,�	$o7�AHm��,kM9Tcc'6*�V��Q����LM��u�X���t�p1��x��s���"�Q�k#��� tRI��.5=��D���"*�G���n�ϣ�DC2���WR�k%R9A"��w��

&TM�0���kZ�g�#Cm0<ZJ9�䢳�j� �:1����;���n��GJ톌�hS�	A��/�(i!Ԭj
Ʒ�XQ�n��y������\	�"rҐ�����U�l�@@�耔?�U���$�����?뚌K��,��7��#�<Ba�M���c�������	v�j��Bl�����������v%5<b=r�j����ك��3�Ա@�b������inQ"a#נ�a�$��.\_8b�n0��ē��+� ����"�Y&�
V
�n�x�]`��?-�@-b০ޭ௠�h��s�&Ip�?MP�YU��_�U�>�D�W�'�^[͸��J�7�� �\B�!�����48�9��̥�F�:f	t��vZ�]�o��q�a
������՚ax2����԰n}X���Y��^�A���&5�M�
�X�O=^5��ضN���*W� e�����4u��Ll����F����n�i���h������0[H�]	?G����@.j�Ttàı�+d��rO��� �c�-��OF�+�T��ϣ�9X�
3��Թ6J�軱�i&C�G�Eώݘ��g��I��\J+(�z5l�s¹3q���2S�b����ҹ;\���F5�:oF���&��0��!rWf��5��Ħ+J3� "�{��P���r�|�Ⱥ��B���yz��%���LF���o�`��M�T͢DE�zp%�
x��[~����$��i\f��1�ǖ!B+!|��_�(-��.a�O�~҂I'��Q+gWF[�ȉ8h���~��{��;-���9=ul���W��N�v+�>�z���*�R9AZ�=��x�'����*{�[��k�䷴�� �bu!sZUC-�a��g:p�:�+T������=�Q�v�B��@�S�t��R�ڄF��^橜�e(��݂)��1�����t׮qiΟUmڷX���=�Nz�$H�9t���1X�B�X>�P}�?��d\��	ʎy��xZA���1M�%��U)�ک�[�U섎�@gB�Y(d�7}�����[Hn��lPQ��2vvĘx��&�i��{+�X�"�'�����=2
�i�`�U,b�gf����G�l��"�#����xI�;��鈸��A�,5;@F����*�P�m��&���������V�k~��K�- ��p���x�n:�>t)� x��M3�)�M�l8�-����KG����8�`UI?���`s�F�p�2�}Z�����O�Kc�f�
�!pӪD%���׷�H�
�8}�Q/�`��>z;C���49fjEPo���X�Dr��;�5���^�[� A67�>X�R�ny�7i<��PI˞S��xMx��n�X�_��O4�d׽�0[Pr�eT��⽬�k3<nvGV�P�^.�/{5^�r[f̉�6�y��y��E�YE�G���*���Ur��%���`��Y
�Ʃ�@�����F1n5�}�z]��<.�W��D,J�d銛a݇�Toud���:D��Y�$��6�+i*$�C��`�S�ws�c'�]!L����qZ0<��Ȃ�u�Nw<�����D��Uo9�i��ş"R�!��,;�6�\(Ճ>�X�>�"\祫=�Ǿ2���`����_i��S̹�1� :#��j\�����[�'��f���ن�V㴴"veў135=���	����ɧ��� M��`���c�5|J��i���'E�)27�J�㯐$b�)��B&)U!���f��A�m�4�!b͆�qi��}�����J��9O���n�8��
�tF^PG���x�\�x�[c�v�RP"?SJы"��q�r����$��Y�l�(�-�P�J1��^	CM}h�T0��	�P�Cj]�P���C}a&��l���Rگh�����@H�.ޮ<ֹuSC�˻Y��h�Ш��R���.���=�C�X�;�J%V�ik�W���z�m�z1$ވФF^�7^�'ۂ�1����j�B�tJ`q~g!t )c!�B��|�-�k!�Q��O\�'��72L+�|��[9�VX�7ڤ]<e?K/��@/W�Z ���d_-Du?Z�s�S2�&:�#�$������tJCe��U��M��;��F��x�jdwv��ѐ�8��7�
�����1��9�-����"ɅR���48k�nն-��\d�p�=��zd)�hk����ۧ��+ �mT�v>�w�t��7=z�ʁ� H3���F�K�#L����@l�[Q�����6�2d<���'D�T�F���-mV+�#�&��0K�R���k	׬��P[f�_AnWL�ˑ�U*�u����$�zfz��F�Ah���B�Ǌ7x����ݰ"�ne��u5�B<7�++�����20ŎW�6�<����ܑuk�����\�@�B�)+���k���M���J�\KFg�"T�"�E� h%�#�T�  ����x�B�,\�b(g;���}]�@~ݍa��V���$��]�+9��FM.I���7��3Lp�e��sfn϶���bs�+������X�4�y��� ������8�����"�$�	f��ri�3������MǗ�W*����P��'R�t"V>�!H��.�҃e��8���ܳs1�� �뚋��k�6'}b̧���3�!.ko/DK�[Q#g7��e�
�E	�zzh~�p��7LP���-fv4��?�L������5��zw������Lӂv�~�F�:xe�~��;R�r��|<7Dת.c�~(r�h�r.� 1O�$� 3u�fj����(3m����N�>�l�|o�)]!�K�r��?�F�ڋM�~��u�������K�$��8A���F�ۂB����E����z���%:|���Tcnt�Ve��=�)[�p(���O>2�W���u�m��Nt�>>H����_C
�k�S������I�/��l�4B(������Q�lcNx���#S6A�s�d�m��6j�-�-,�C�7�Mr�x�61/x ��QPR�L�㱥��;�m��(=���
�#���ǥ%Q>���/|��O�,����F����\T��L���k~j���@�����u�.�"	������G���Qͭ��a��:��e���>�6���m�NU�1���a/�����d�-�p�ȟ�t$*x�hgl���{X��[7#�3K�*�~��Y��RN�7*+�	���J����L�������Ȏ�rO>x"�.[M_�	_���/��SD3���/�K�+Q)�РK]���ճʈ� S�K�gf�܀+�D�k�y8x���o@ݬ�	(����|�#� w�8
l>��������3
���f&����Z)�ϲ�"a��V�����' �=��e c�8����]������0�O�h��y�"�������W3M�A��\0)k�ET3�q�0���>ҳ�=FY~>�����:9�_t] �;�ne��O��/�X��R: ����uЛ�Б��ۨ
��na��y�&�{�RO�]��p�>��[
�R>�����I�d:�H�N�1�ż��՚ghM��h��_""���<��lHaoh�/RW�;%��Q���g�J�r�
�F6�1�9x�m�����+���0ww	��������5��;!�����n�/�n�{ﮮj�v�gG���z��y�?(訩P]�Se�[�P�x����8�>��R
e��c^MI��T���7�#�ʌt4���h�#U��NKv%�9L�U�.��9�U����6��V�B\�ِ��H��b��}����"y)��tϢ����m�[��^L~ng�p���;D��|�fYg�՚�Z; -<O2.���{�;�� >���Sr�$f�X�db�ߧ��sP4�AF(8EH�v�ӧ�%��&T*T�u㋐R�tI�=�����U�|L�f��]xL�.mL){Bh���$�-)�{���ǩ�M�++�M��d��G��ik����@%߬5B���Tk��#l��$
y��f� �����*~�~	�h�*=Y��fܢٴg���ǐy�Cذ�	gT�F������~*gC 54�C�/��$6���y3�^yG���>L��C_���W#2�#���8"�V����z��hm&7��sD����T� �e��Js�@��OC�ov�$t�)� ��*�@�Xտ�$�����%�Ù	`<g,Ql,�����S�2h�U�|���e��Z2]C;���s��N�7ҕc�~�Q:B�$C[���F�dn@L����X��/��;i����%��~l�*���L�G����k�
ޕ�F'�)�1cD�9'Ș���f$���F��ؤ�W�_�c�>oz�$񾅴�E��0�����*�7Su���G�]��3(�U
��'�@x�*-�^чY�ʎg�!�Rѹ|gCĞ8�̈ޣA�
����o�J�%�)~�R�x�%I/��̷�I1C<��20�kg��Ӵ�l��i�d��CM�3�_�D�<�|e��O�kII�_%�j�^7���L��ߐ7�T����B�є�D�C�|�`(����e�B��8�-���F�G>��2�E�	���K���C
�t���$C��;�5�uQ�!.rX�W}�҃�YU��8ԳZ�&�{��ږ��x�v�Nɬ�;S@�G�P���%���d���x�|g�}�t�a�OWC!�R���~V+�P����o�HkbX-\5��՘�H4�%e񵓥����~�����/nO�[f9�n���	�,	�x��r��Qgְ	�(�pH��$�5n�>(�}��'7Ϭ�{q~�솳Xı���!�\�����.$h>� X��S;ђ�o�~����a:��c��pzT��榳����\|U0L;���L�pK��%���s��.���v:k6�ٱ�R���T���3���Lsь���K�o�9�����s7�\~�C�f�*�h"m�QQFK1����V�u�0�,�#��Nvc}���xC�9P��C�_8����^�&<`L��E5�ٽ}�޾%�_zJ��dP�7��C�U{s�SP� -�e�l�hG��p�T-�Q��:��tw��d�f��j�\�"L�����'�е�d�з���J�P�B-�Y�Uh~-�� ?nrN\���8�u3�7�z�^jԷ?�_i�uJ�~ū�)�����nL�]����`�:`��|�թ��+�l����+��k��'�R�h.��;���**#�0��,�D���78�)��%F���EV�*����C5@����P]s���	I��Q���o�i!=�A3p�h��I���
e�߰R�y�oR���KF�^R���1�����y���� ۛ�I�(Π�W���8�#m)K����ۃ���x���=-������nS�8��ܟZ�&�D��4{d����;:?d�T��z�����k��I��Z�����an:��ԌP�����7�g�c�fE�5�[���M#G��D�<U�����S��0D��ԁw��+TDi���)6;CF��5y&Fzc	2�sr1R�p&�����鮆R60��T��s��\����|�~��������U��cs�ϝ�>]��ރ=.�i�g	���n�x_���BI�L���IoƔ�C�^������RVDY���ܞ�����5�^�
ˏT�|��5��T
�Ԃ���TTV��t�G�)���6>e�|g���	I8�Fm���S���^[�n2@��ݎ���R/O�+$��nn�-�@,	�����}���`n���4F߅Rw�� |�� ���X%�R~�T%nLO6	��4�df�w��[��,!�[Du��UŬn��!-�����u�N��ςz�m��\9����wh�`i���,�Ҁ[jz�3h�rLJ�0vۄ����[h�+��FE��}A{Rp;����~f<t��	��Qmk�Ty��	����ַ=��AcB�%�#�c�8
��?�m�v�	�N�VT�3��C��}��Yẜ} 
��(J 0�C$�V��+	\�w�%�'T����l<��m��G�#�Y�.#>a�X5��q$��E�����D���`�{+�#,��:yi�8�=)��嬿V޺~��m�������:b�E�$�*�Hۆw�Z)�n��t��� �p�!��q�B�"��椴�X�Bx/Sx#��4x���4������*�ɟ�`@;�$� �zU��M�(rtd
��u}��d��/�J�3Oy��T��s����l>|p*䣆j2E����"p�N$��H\h��F��?֯,ܘ��P���+R��*w�P%��o�I�i,׎��a�ƫ�������$	�����.�RǦ���>���,�D҄&���G��k���w #�
á|�6�µ� |R�._@ _�FV�>>W#/������_B>n�S���J*fk$p���|�K�j(��8�Xǖa�x��q��eG1}�3
�//I�:;��	\����8Zr�����rE/�t!@fu �^������?-�q�I�F��s
[~�����CS,&�����&�0fp���ٯz��H������=o�;��vgUř�WĂh�@�5q޻�0j�d`�O���ձu1����e�y��!��dZ��`~Ÿ����C'�MR�t`��#h�#.G����v����*?/�����^�
�N�^8��O�2������&��6d ��w�m�LK�c����pS��Z�ڨՌ+KP�`p���=�ТY ���1W��9V��?\�����\�R�\�V�s���-��av:}�*�����[�s9����EQ֏>�/�	?��f�̻[��	�!%MW��xm�d"�Q�SJ��� i(�A��~�Oo���#s�&A���|�ЁDϥs0>}��r!�*��D4˗5(W��|��W>�G�ợ4��f4/��e�s��l�I��H���]�t,ymo�~Տ�Nr��t�=�Z`n8�4���k�L��Y����������{vN8?�0�z"�G�W���`<����5���>�,.��(d[3B�:K �;E���`C��hO��,�$�J��"%���X��q��"�.v1���iP���Oc|�C���.�+�m�c��|ٰ`k��ƈ�k$�� tC�e6|nի��4L�'>�t�e�-�$z~���;���+�ֽ��Rm���ZZ�w ���JM`��&�Q��h@�U)%���yj��0�G��n��eo�~��m qE;C�;# ���/���B=�,"�
'@�%��G@{���:�J�:7��E��=���Ly��s�ߏ��\!�~sv����F@"թ���5���"�I�|����n)�&�ϡ���s��9Tb��OPվ�s��"s^�5�%�A����D��p�FY��O���Ѱ2�rI���h>������s���]o�TR�߽�u��z��������t���"��ڱ����?�p�a�fT���=�r�&Y�ݑ!����S�G���bw���k���(o��x
�d<�+&m�D�"�ȰPK�{��p��ѡ��M��S@�q}�=h�ׄ�y>L�����깴u����A*W����0K�M?�/ j��m��{T���>xVf}m���rh���\��\�U��pl�XE.�l�H6�Js_����>������8���iX6 -z�˴��n����MH7b�����7[8��M���K"�`����d is0I�hQ-����,؋�Z�:c�ݛbqk� ��{�|�����e�������M.s�����	��3�ϥ�� 	hW��9с ��k�=�|8����ȡ�X���Ĉ�s��wmQ�&R���[�^t��7��m�%�u>-iӌ��V?�`�����c���ܴ��x���OtZ�@n6ȁ��o���ra$����\|���)���s@����)����/�$�3�*	��f�9��uz��
����n(WG
0Fj}��[@<&���q��lq�L��[{I	�ޝ+���w<�����KK�Ʌʱ�ރ����E�7�ű�&	���%��-lHZ<����t������PX�mݤ�����d$D}K��5�%�+�L����Wk��mG� ���]�)��G������m��n6�L�f��[IX�}T	�]Hl��(S�����:=gư��I��۸�N�'��]�!e�pG=��Iq]����C��bܓ��U�����2����+m��{�`jq�h�FYv��Ajn.|��B�"0^�.�!;�<)��\3ˀ���.Kjr"�gCu�md;]i4m�?!/�ܾ�$��N7�X��1���CDOBM�8k�A�e2-6k��&�{˓��Om��My�ywvv�����H�|�)��TgF%�'��=k��=��ïA�`�KQ�ZT7q\2vk��U[�!��7O?��]"��a�n-��:�#R��������)�x0�3_f��
�D
��a��NoM����wx^���S1� �߲�.9��_��MK�v�aJ�x��d�
�,Y�X�ȫ��N�=�]�7E�3�E�l}J\MCV�#�b�>��=�CM7���c���t��A#/3W
����M0�[VP.�{����9�� ���Ck�O���h������OvEߘ�̷��&�I����E4WcY+���s��.7]>t<N@ J���g�z���Fce���)||�.��Q�5�,��*��$�C�v�Z 範g��d�ໂ�z�-Ԯ�#�a�T,�h�[�*K�P=��C<o����u��B,��	�N�����k��6�z8z�y�L�ʏ��ټ��S��('u������hؓJ�oع�ȅ!ӑ$�O��JM��P��!�Y3��Ƚ�3����ɟ{�,9�{��Z�����������d���:�Rˠ��%�e�bg��uD\𖾇��gf��8���
�[qI��d؜�P�.����4'H��P.�Q%|t?��"�w;��Ҽ5�D�l�&�Sh�J��Q��F��~L?�ȉm�s!�A��Z)�޹E��{ۇ�G���8������{���J�� ���E�#�������Rb+�4`L6�G�|��F�K?��r�g��IWйH^�q-Mn�s=u�۔�d���3�&P)�t����O������x����I�g%~6���Y=������5�9z1>b��O�G�w?Q�|�LP��l��U֢|��#Tc#N:#C�|�v�\>>�Dk�W_7�&P�+����^�>y�ݳ���W'�Dfh@5�³mнVe����[K��B�6���]���u�JJ�B�:9e�q7����/��3*�r���8��B�GjwP�G�U�)��ſ,��:W�;��qaݩ8`�������%WQp�])���Hʼ���G:� ���ViN��S�D+��b�6�?�a���3?]*�r>h��<��������݁nX��"r�*���Ɩ��˕|� Z�A o:�?�x����>2�~���l�#ξ3y(��3�V��� �Ԣ�
���7�Ᏹ̙8��L����徾��q�U�s>�p-�٥{,�˔x��g�Z���]բ���/���,���՝���qsu��`BHþ����5�[�ԅ�������|�A$�a6�$fB���Q���5�x;�F��G���c�B�
��6";ĺ���
��oW/h�3�x�K`����\c�Bם�ul�s�)﫠et���[�U䌄������&�܌n̯g���(`�E��rqqI%ѵ�n��G��$p������Ͷԩ�\ �e���R74990�؂;�+ֺ�����W�3h��էBO;/Jb��<��������[�j���刍3�cM���B���⺫�Z�|�s�7��}�[���Sjf!���sy��`\X�ɾ�~^�k�VeI;5�=R%���V �g�#Tk���C/��i��!KL6����ˤ�h-�)cv�5�g�QB9uz�>�0D4к������U����u�aA�ns�KE���Y-���:P�I];�����@���/t�=.�r�6�ʧlj/}�'_1�
���P��7� ���S�l�����r���$!d��tpXr"�Z]�]��^N�(@���9��t[�Qvz@��fD|���$����Q��{`Ne��k^l���`YJ�=s�%oqg����������៾��;��^s��ȥϴL;�e1L��(�1|��{���w9!n'h��'�]3h�]���
�
:NЋ������|�A��wd�(��T9�c�s��*�M�sd�����7�To�a�.Au���H�gZ <]��ĭqǍ���C+����廁ҷ?�ڪ���&�bp�)~��2�/ʸ��45�e�Ҩe�h����3߹�<O�`�F��ߑU��0Կ�z�q�I�ND��w�xq����PP4�d�n�]�<,���xI�:)I�ވt�|�o�7P��?H���cסMA�t%C*U&�m�����J�i�ONI���9�%�S�����y�H�֮v�IU����bEq'��<�"CKh�,��IM�<��NȆ�h1@p�8�D��t& tlg=<�X��ИKԡC��;���{p��!����Gڎ�������o������3��j+B�����۰�f3snbxU�|����3p���}�
ɓ%�I��n�N������M�&�8�ZP��eԸeذylKM��.B�"@���*'��M�
��=�CR��&�C��CY��5��M�n�
�.}� T�<!��s��(�G�f8�+���S�'e~���$�-j�yk4}s(�
��F�:���{�!ʫ+�D*6g����PTs1�5��l�uR�&O������d5�9�И�=rũɱg�)B���ir�{8#q�����3CX�{�f��M%�x`�'�BP� �K���lI�����9����_���9� SG�;���0O�<�z>�f� �]������D
�f+�����wEy�ǔ���-��'0��w���,�ʌ޿1�ډ�� ��d�	L��䧘],��|�'P����S)Q�;mTq�О�H��.�Y������Y�/�������� òu���j�b!P�4,�6c<ܩIs�6����x�ݹ1��ڎ��J�,� ��%���18t��E�&l�4<E����F�[�5^ٟmvf�2��˷p� � ���<��P靯���˸dG�>\w,�F������W�^E���Jx;��=���/&u�7u��r���A���|���ɼ�0��1���r4<�w����ƪ���YE����z��S}HYY �҈T��Z���/�:�E̰qI����:���h��;��OƗi��Y9t�w_ �|U����x�]�;�Q��<�?��<a�C�-����Ҟ���E�X�|Ę�{�rL����ƽ�����'��$v�I���l%!JU��G,F.�"�|P��i7<���G91�����-|Q��:�W����)`��2��ǔ������^�t�O+�X���xzY��1ҋ$�|ْ|�>3m��0����/��^��6	�(��V6A����z���������g�v0xY�X8
Z$X���t���Di�1�.�2�[ק�ݧlT��\���G;�s$ǋ�S	Q��2��H�	���Y΢e��}W=U�ߓĹ�	�oN4+��=Ĕ��}�Y��J�T궴%�3���x��t���]�27OQ�>�*�7�`0)ǽ���Jo:s���K��@��W�f�x��y�z90$�����ǿ�Ym�Z
e~�§�$�l$��\�
�lb�o-�l;w]>D�a&iMM��r�^�l^�	N���>.5�|H��o�.�� ѥ�}*����.������ɚ���-�o�]��&6�`�1��-��P]��k��.s�������P<�
���~��:O�6������.�<���?8�@W��@dg���n�F�{vl�b�d(�6l[�h}�8#�O@K��� e�'���$����-��M�(nv�b�"���R�[�~���gCSQ�Qsr��� QpL�S*H"�5�g�)����~����wlHO0�1�yZ��"F���@�'�o��9�]�o��Ij<�@?�Xyd�A�z�HF����C�����V�"�tч�ͬ���)s�n�g��6@9���}����1��	(�-] /�Nk
��߯n�?�!��8QL���\�dG��xx�z;��L{��aS$���|�2_֛޽��N_��/��5�o|=^7iz�8_1����f� w�#4��x39���z�)a�ڿ�$�t��wH��ƈ�7*�V�(�.Nn����Q���b[���ӿ�w"��.�vP�w���]���2� �v���\�V-*,e�=���]�s� ��8��;�#|�fߢ��t��;N[�C�ݐ�ܠ0?`�Ƌ0�wQ����"�M�<K~ޝ�}��"kn:�*-�'�����Z��5�����/���;�S��u�v\�my�!h���H�Ò?S��m��
1�����-%��v��>���0������q��֖0�Y�X.��f�{���N�%�@���"0n��_��$�V7�>��&����u3P�&�w9�I9�{�c\>�s��4O�·C��W��Fe�U!�V����Ȫ�av���GHN��T~�����g�����R��V��� ﯚN֝�v�7�</�=#�!$�[X���?�����ޘ�<`CJ��ú#�31Z�nD4�a���1�����*h�>^O��כ���K��^�V~�;�0�c 1`�w�Phi�%԰�V絹풦�����K��E�1�H�����W���nHJFUTk����0t}�Jn�EѸ�U��)�M4>�x@{` g4��%��xC����R��R��d!�t��c��d��["ᷱ�HK�޴ o�KM�uqK�� ������b��)�5��f{yK�b�K�g�j�����^��A�c��ȍ�C� H@���F���jѡ�VԀ��R���_����]�U�l��)��������dN�|���C�?�+G��9�W��61�jn�����V1�Z�G�ձ���hE	>C�ӫ�e2N���rw�o��s�RVQO���z�'w�]���Bk�{�?��=�Q=;����?��(Д7]n=H%�9ONϒ2��a�� �b� ��8Zi�p��^�v����#m�8�E.m)�Q�b2g��~S����>��evp�A_Z����r)Ó�?3z6�me���O��z��xn0|�*dE߇����0�r_��%�z<����#u!�~�;ۜ^�JF��X�"ҩ�v��ޣda��]��l����8t���F"�V�Zl�M;C&�9���{E���O��vjs����2L � ��7�v<��>��e��������9ݥ��+q&\�����V���7r�%�-�ѥ����ԉ��X�i���?Ü��.K�����J���ѯ\�Z4U���l�$P ֳ��O�O2�#�r9۬f�6��;>�xH=j�DR�)�h}MZ��C^�u�k�8��,l�����;Sߌ�����{�䟋EK�,�[	OSaGN_������TR�����S�@��6��Ow{��
��<�%c�<ޕ��|M;p#Ƥb���#�V� �,����+L�P嫯s��k��1a=,�JNcP>]��\'�.�A1J��u,���������/ˊ��q���o�.*/�co��[�Y�R��-�&�Vq�*h8�dcW����#Y��tX�ۂ�Jo�z��=�0�e
*&�S!�q�����$������k��4=|_��8T�c»����a䤒[W��Th=�}��;a�U$򡚘~N�HtRi�6m��ᬽ^c�z5g'?&f閑�OV���1�� 4mZ�+�2z%#B�BE���%��l���i��6�Iy�"�p!�W�b�J��Sܗ����ܶ6��݄f�i&��aõ��z_Hｰuzz'��k��6�9O�P�t��r%�Qd�|ƒAp����>�M���h��։B T�d�F���{|e�0f�$a��{�i)Rk��R�O�<wsYuC�IY�5P��34E�%X��#��9���^	�a
,s��b(�j%%�:��t���M�e���ݸ���qȕf�
�q�E�銘��~8���c#RcZ����QS1�YC�������W�8l҄gPxD����P2�6�+��voV)Wv�e��6a� �c���ܸ�b�]ƶ��U�þI,��>{{\ӟ�Ԯ¹��1)������oM�g��s�Jn�����^_mE���\L���D�G��s�wQz��8?:����`k��tu�8=!J�
��� b��3���KG��L	�8�z� �PK�t�lC>x�Ɛ�F^j������=�>d�z�B�S�0'�nm�2�+IU�a(�3�|��ͻ%֙�1qj�ƩW=Q�Zҋ%�A���:� p�]�;�v�}	�&��>���u��z��Ֆ{-���醦���Ax��U��_Ȅ\'�V��bu9�w	�Ab�u	�5�SzFT.�Ԅ~s5��l�O��o������,T%��$�Օķ���HA��;l�n����n�(hy3b��q��ﷻ�4���~G��2������ۑC��� �XR��	OC0�/nC$�I��^B��Bp���x1�JBe�So���Nqr 6��>!	O|�|�8����gN cy�<��D��J&�,B�D�iH9��3�%���G�61
'�e�T��
t[	S��D��=����8���N<f4���M�OFI5$mGx��{���R7�³k	�gϗ!W%��#��2C�0z�Zi�v�(y��z��/Wd%��@y��i°ȵ�ߔ��d�/:B0���e,$~�k��p�B�]����Q��Y�?����d����p h$���MSq�W�k�E�/`�;��TH쯂�N�����ǿ����S�Jp����+f=_����ݴ�Fzѝo�������:�)E��LN�&֌��{�n�1��M}����@��*1TƎ�,%���֍�]G?�|��1�p�z�9:��+J�b�Ӗ����G�Jv�f~�I����ټ$�v~ڿ,�"��mjs�����*_��N:��d�1�#?=|{�ڽu�9��e(��A�p����*�ۨ�����a�jv�Q;�.��7�B:�*h�mkO8�)�q��4�r�W����i8 @�	���\���{��yA��M˦�jDz�������1ʿq���=0�A�%%����BkU�����1�B@8z���@ԫQ?]MF��x���),x4�,+s��v�d}��G:�����@?�a/�~-W�OaW����s�����ϳ��$�:���o���h��9����g��&�Na����ho�� �ll�s���	�NO�p*mw�|Q|���`�� ���?z3+G5b�+6`W���y���
h>­N8>K�xJ�yQ`d��#<9�<��,��~��$/�f�b��Ts�P��^_�t�?��R�R�9�VB_�~?'G�(�s��X x��*�v�k�N�>$�[�pQ͚�D���ݪ�
�w�����܈	����품;��]h����N�2R��E^�������'�z�ffL�b��4�k��	�{}���G�rI���"O�lr��]�;��?8<;vߵ�
�Z{�og�˸G� Ѧ��V4���p�y�Ș��_���%����D��������{��2�5��{c=7��u��?9�F���J~8#�4TZ��z��)"x����_%!������aA�*��|"���
8"!��Jv�_�D��t��0���ņ�KК�1�֙z�A\�K�}�7�y��6����@Q�;T2�e��fM�	}7Y	U��UI���� *������BY��`,�L �ɇ&��i�}�e� ciu*!�\D�wԀP܀PT�6��1�'�5S!��x�,�gF"FiL���j<�|>��������N�q�-[^�&]&?R&�&R��N>ܐe܀�m�j~+�W��T�������+C�i3���;���>EقL�}K���p:��.
��K8g~���3�\=�����c��B}�$�5w3�9a���jOtc��p��P���
��s�p?�x�H��$t����k����TB�,��_2:��v�<נ�<��K�q3�見��2S�5H�����ʊzB�`M���v�F��z-�*����zl�u�=�HZM�Y�sc�����%�w]că�pb��D��s0D��`_�����{��W&X�y��n�
pdܑ�me���ٺ�R��Q󦉃��v�D2{xtq�u�L�I:�M�4�ޘ���A:�md=�s��s��Y�Y(nv*�<;��툚y�:T/U>ji����<�\��H>R`T3!��w�!�����d�Eb`dd��V���1f3����JJ������	���D6x����M�eVs''�b7�%��B]&铵$��6�ɓ���� :˺��V%=��)$8�5c��.:paϏ�6�K��:v�GgD��ms��;��|^����>õ^���6^����(�6�������=�������������j�g:�~ȊyDpkӃO�[�]�=X�r`�\��y["�m��zٞ�Y~�s�=�����-,AfTV��ʬx� ��V�5�����\�y~<�!$z)M$���w�hs?:J�h¶c��_LWߒk>�#���ri�<=/�:��OIM���T9O���׼�ZJa�NIH���o��r �}���xy�+�bEDDL�*ۣ�CC�cKɦB_�3�!��m�@6�n%��O*U��U^i)�e�������
�����w�.��HC�%�\�R��!�J]��XZjr*U��&���DK�k����^T'�ν��D.�k^�� �ũ����P�̭s����-��m'-�Eh��JE���B��㢊�G`��;gp������2H&0Pddd$O��\�`��g��[;=���a��]�X��B6f�ɕ�X9�,���B�e�R�]�.��������s�S}��h��#�C����འ�9�������n^^N�A��FT�k�?	���9|���Pbfw�p��4)x�����=��RP��(|Eظ�>%/kf����f,c��J�/����x�D�������l�#��2 ����=V����L�^����\�zNGG<�/�G<�xK9�ŏմ(�Ϣ��ClQ,���n���d.�`��ś�eai��Eް������s�3�=㯵b! �FU�Qn),@ӛ�\�sЍ�턌~�̑ܘ��SnC%���ŋ��j�v�:�`��$�U��-`hE`d<F}��X�y�hEc-hlą�8:9	ݼ��,=H%����z���|A�����!Q}�"A#$$��T{�l�a�jJj�F�`f�4i/$=��2�.P�Q!�e��E�z�No�Ҏ��Az@#Q��T��Ն��]`s+�8;-n�tum#$-^��m����>�ñ��.-�D�����	A}�HFs�!+�?P���K[�����򁶡���#s�1:X�����*���t�v��8[���!��3W����*^�k�V�h�:N�lw7u���oʎʞ5Y�ª;*��3E���- B���{�rmd���8����ZNl�t����;��Qҕ���d�B��$�b��!"� G���g�4~��2� �o�����\_qP_��[���^����HD0�U� P�1�>E����M�i�<�azT�����������Zo��:��;�!������e+	���[\��'[��R��ѱgg
���RRd�^�=�Dǔ۳S^��d��g̦�yV���������z�I*���8?F�)��c�Ϫ��� z�|߇���?�ump��8�r"!�p�ڊ&�Q!�wA]�{}�lm��:�6w���_Z�!��[>#��bʕ��c��Y��,.v[PQ �< | ����Bx��:_�Eb����S��B���l�jɭ���ҹE_����r3)�y�����]��N^�����ӈ��Ě�<%+��9���p>���������|��q��Mi,';щ������I^�'�^-'9"�	=JB�F�J#g(��d��Jr�mw�q~:�\��[�~u��Dӥ��y�0
R������Q�CsTf�^�(=+;��k^3�(�|5�S��,�^�Xx�};K�j�m]�mr���c5'�\m'A����P!����IE#��zv���=��[����$��������O.�^��Q$��J��^��	�_Z�>����U�)�(en̭��5��ڭE���4/9B���&X�˫�
qj9p���	xqo��At,���ˇ��:)=)��\:*�f�%9a��.֗<��rF��0��h_+J!;\��j!���1�t�����*!:A����!���h{z>���B���K쀱~2��c���wv���s���0^�%J��🜞^�_�u��U�hh���cH�~Wd���[I[Z�jؼ�������J��^��c��R~n\'$̯���!H�P��K]��C��'���Qo�ʁ�wfԬ�k����zRZ��9��_�?:"`�s���~�:GU �uѦ1�,_	H��j�,�����&��[��,�w:����aja��14�/��	�!���l_�^J��q�S�Ǐ���\E�#�F�-כT4ur��8�I��$W8�,�Ȟ��M��;ie��n&�6G��r��e/�/��:�t�T���Q5�5�P;4�sY��9��:��\��{|_s��~�5E��i�C%
�6vv�������R�T�MM��R\<<;p� Xؙ�ZYx�Ύ�ͨ��NB��n���&XBŝ��T*��ݢ�C��,U'��Tԅ�<�>��(t&����B�֢IJ8R4APY�� 6�����N���3�������"_M�-�v�1~�ų�B�{^5lҫUG���7}4�&e#�y�$�%�l�bC��A�I��6R�Oc�0Y1}�#�^�0��6����}>��|�   �YK+jaa!K�G9�i�����X��8O
?l������O����G=���|S����+�y�{��ḙ���T��O�[�kW�b7���<M������o��&��q tP����{4%`��s�W�"��Y��O�z�"�ݙB⿎γ]Z:c�o;�f]맏���!���޶���|�quh��z�[$x{�)��l�
ժ>]L�<��:x0����x����Ύ�[F_���,x�qp2�����Ip���W[~����[5�j�����J��YEv�a7���4%�R=n�F��s��/�#0�^9+[�ޔx����"TT[#�Wv��wGQ�E���K���k��ޱ�wV��.���c�z�~6b��΄体��Gk7��)(�Z!=���lͱU K.ujz:ddD������^�1�#<��-[E_LZN��'�D�n��:�_j	�!�Ǩ�w
����\-��ag����c��w�2��שIdX=��͐ֈ�N��x�T�q{[��u�V��mrPw�*Wj�6R���=F4m�7�q�W�G$�S�r#��Y�Ë��b�6������Ȃe�<>x���ł���'�j��e��ں�+�Z�0�͇H����36l�ʹP�K�����K�iψ�
L��'���ž��n+#�ϑ�%�_�t�3[�c]6~]�����|9�Z�	�+蹝�W�)�Ď��v��/����"���.���ໟ��L��p7IT����ʈ����%Ov��h9��x��p�K\�$8�É~(4��:aE�a�l\i����E���ՏO�;˫&��?1�� t��.f���@�vbUr�(��2)������k�1�c�������v>đj��J�y����]FfF��HxK���ܜ���t�:�P��w~�ӎ�T9F�n0�hUo�^N-I��i�x�b�D�`IO�3��) ^��Ak�x�d.�q5��nU�n�p�,'���H��{��Q���ߧ��1�I��Lnk'�\l,פ�0��q���7mH�|='��x~]�n��pt]A��\���3��m6����a2DvW�Y�dD��%���6����w���My_��6X؁�1����P�=����eh�O(	-�4�w"� p�|���.(��M�I9?r��"��EPG�@��I;�ů��� 87P���U�ڡ����=�c�6G�omaҾ^{]M��a��l+�¥�R-���[�$������nO;IC�7F�Z���]B����+���mwwww	��	�]�����ww�<@p��<�=|�����M�95̜3ջw����)������.�qs�I��\Ґ��w���"��h2�f��D�ӹ����=m.0�M��iæjQ�Y�G:)�q�FP�N3i{Y~S�6�z=�/�<�>_i��&2SA�{zu7�%�Z��]�05c��Wx������Q[˜�gFO.rp���r%lY���OG�ɏlg�{̗Ȱ�Q�}��I�0����|�+ɀ�_�̌�kt�"�Sh*�Bg�̣����2)*�F��L�  2�a�&�x���<�E��	����F
��z�Ϟ
O��<�J��9I�蚴l�@2��$�:���)4?tf�#s��rJ*nm�t_O�z�箿^]jhb�t��L�����~���u$�,�o���1���B������y�K��`u�������������s���jⲍ�����ݟ$eӅ*�Ë����-7|||1��6N��D���u��꺰�m=0��l��!�YOmS1�=��"�_r��p6��?�M�S37�������qހ��ɜKa)����Tbggګ2Ш�ÌW�X}�Abw��g"w�K���ۆ;d�E���o��x��e�M:%t��#�!����igm�����a��
�v���q�G��	r�|<[��lc�->I���C-55����8xF�+��?����Q#M��o��n�.v�5٣E}C8��U�T��8w�m��	2,:�[���}l~p�8z�P9��w(�yH;H`�DzTn���|�0����Bg��?Jb����e�˓X�y�`��85��_�p8l� w*��o�Ý�
'�}%]����I�f_L
� t�'��^J��s9��z�ږW����`�||�|�t�!�<�x���G�}z����Y����_?6'W��	�3z� ���%Y|� };,����Q��n�C߱k���Fc�*y����
ی�<7ڟ�����%>[�O�	��3�\�}�?o@�%$;��r3����>=�)[�}L��iZ�@�Sۆ"�#m�Rw�p���nIy����d�1w��
�t5�}�^��{�x������D@h�(f���;����%BNG���$P��h_�M��v~f�9j�y4�R���n�^�W����dK:|\�J��b)NZ��B�yM��v������2X��/�I,+_�i�n����E������6/��W�l�3����A[!��O)�v�h�s@��\a�>^�9/��(�e�H��u; ����|�5 Tq��E��B����
��J#��G
��z���ٟ�
��
�$O��F�-�*����MDjFw�Tm>�9���&>zƟH�0�w��$5��U�S%�C�� *���&��%�x�Vоb���T�X%W^�mj�k�cN����3W��2V�n�j�e����4�������(�Da�)��>�3�@A�s�^j�ұD��#�@���?���ٙ ���+��j.�L�/"��NcB���3���(b�:���.����Y-%̠rMmo�ꅂVߺ}ֆ�:�}��+��\5H:M�������=k�È���O�U�`��C��=� �Z�ky!��?	Ǩ?�[�����o>�;6겴�����:g�S���Q �� ��O����� ��ԸMm�/2����d�o�7�\��X�FI�.�b�Қ��5���&\�Cx������a��bC��L)��t�Z[I��|𶣕�\Ύ�P��iE>O]��!i�)��Ww��C��؉ �*F�h�?Z�]�ag'��m�V�#�3x�b��,E`歛<�(5���k@)�.�QqL�k_[��ɺ]�!>�)AV�X�k���r�HZEΎa$i|y�V�ى!�"Ob�V�>����mӣ
|�uj{A�Ϸ~"6���N-���m�c�G�����ⅹ9��B��r%z�D�����׏@y�K�(�;�5��Z����vϵ�`���r�AyU;~T!��`�ϑ\��!7���=�(Rk/T�%2�<lP}z�Ap�j��b�H����
��8��3��oM4�e̳�Ą�Uc��p�V������{�5����0�Nj��m9&.E�1��T��kyNk������'�z��#$�n��6�N����-�!F�󚠮iHV����e�,
���5un�y�L���cӝ����EJ�b����kZ<��w�"�˅��k�m]E�:�t�j���1ouF��A��r5MM8�?�$�LHX�5c"� ��M�&���X��Ҡ�|b��<��۟��fP�tx��S]���o���k}��Bh����'3�-������@+헝�e���M� �u%}������\���'c<���O.�x��!f���(�w�� u�}c��G27�IS��Uw��+��=t���A�,������	�W�����G�q�Ӌ�p�c�i0Q�O��]��о�T� ��md�\3���s����(�9m5��>IXd����Y���d�F����S.1o� $��|'�������w�Fi�H;�(��y�����%���������f���*��e&$���fވ�_�� x����Җ(��PNww��v]��s�\'777��,�zk) �	;��i�;�
��Ѡ�%N��J�}�v5�� �GRpxh���4���Y�H�]j����\vдXxt�h�Oe��Vs��q�?AN{k��iq�����+4nS��Y��ڶ�^��Rl�'�Dj
�8���?�X\I_>)����*}��K���}E�_;ֲݟ�N�|�u�w��v����i�Ae�n�,�_[�MY� ��*]���0����F�OvN�Xh͒"G�v#�z}�K����M}�x�:���:\�LޗF��g
��&�v��4ȣxq�p��s7���թ�����6��-�/^����o�d"H�}���0=/�ϊ�����[ ����o��?W$�/��O���qV�51�U��Cp[Gp�ى������A��=QB �غ��> B7����'�U�n=W����??�!�0)�ݸ5@�wY9!x�0l���1:H��l,�H��� �J�hn��~��������cn �O��M�4�3��5b��5�)2~,�	��`{�8��Jk"7��R:V;t�JW���B/�1?Km`Ѣ"�I���]��@R��g�S��۔����GE-�W�L4�z�%���z�����C$�Q��mthk�ed�[<�����4M:���H��7������(W�S������j��T%76J	:��"R��k3>}�e<u;�@C�eGG��3�;�ܖ��0����aa�Ez]A��ᛔܐ�r��%����TW�|
Re4�q���q@pl�e�͊Zs:ކ�u�!l� �N͎��FK�U�KIO�!���>�$R��gȺ�KL�tB��-+���^p-�&Rr��c����b
�[�X۶v?{���Ģ��,S��y�8)�u��	�v$�R�����<m�zs8QB��e�8�ę�p?hN���#!{�������&7%���zE,h�0�W��}�?�����.8��.�5h���3��C�C�ο�������z�ɩ"�k�f�2�!醾!=O���EШ�Q�Q���n?4�|�~գ����Y�r�C�~�]ÎF�{/�' ��.����-x��3���H1���}�_@��E���yqИ��+p�%��!ʏ�ի��}4��ݯ�W��>U ��)��v�o�z>c�U�W㑵��>]94�@��	�b�z���E���F��,��	�	�����I���T�8����`�?���/* �p�7B%�
D|t�&��In����ې��!r����{!!{�!x�4L�z��^�||��*�rz��E<ډ�7�Qz���.:
�<�ZZR"�����̃�O������ϳ�	絭nq֫?k՗>�c`<�M_K�^��'��vXwn_�d@�e筪��ϻ]���[m_ݞ���<�QH��9v�+�vW�����j�p�
@b߄|�A	��n�����f��2����@6����2)"ER�xe���;�j��s�|�Szs�C+��)��M���QZbk���(b&d�r��f�e|_������U4+x	�\X�W��X�"�.v�I��q٢����~�B./a�jp3M\���7�>�,4��teJ^�)��F~�7�5:)�4ut��D�#A��UU���F��!p�Yb����q-_�d^��
�	�p�T���sh?���`��tp1Po脚E���}�R6�SCL��1�J:Kt#O�~�[���E�ɠ�c5��2P����e������,�ාb߹�閭7sQ��!��Il�9b���A���*��GC$Ⲛ��� Bm���.H�P1RsZ0�b��o�J�@�)T{F��|��#��u�	ߣC��`�=�<��گ����6�򕶤D�^*�^y[|l��7>�͸���H���87�1�gd/����E�i�_6y����R�.��b���T�_Bp�4P�#Uf%$�r��aGbU�%!F�UoH�R����W�{K��8VX�VDL("Pn��ku�k�sǷ��Ya��m������BK|�Z���Y뱬(X���bnb�,�{Ǧ��ο�� �d�I)n°>�46�agt)��ށ�N�~�ƫr�Q/wJZ���}��W1�hѥ��EP�2kYfp�o�����^aQt�
<�U�	_�$%0�6�K��O|��Hγ��ư���n7X���I��Ƽ+�'	0�4~3��3K��j_�n2]�����e(��`"�s3�x��O��>�}���FU%�
¼�4�MT�e��䏇���q�9��*i���6����w�p�'3�Ψ1��N �P�g��lK}�F�����;  �K��	b��2���8D�c9��z�d<������?66v^{��U_�PbZ�v(^�*2e9#�h��Cgu=G�4:�x9�A�٧����ʋ�y�6�7Nz��B������q/
OF��>�B�%~�^��<�Y�=�|�~��E=9��r5.�@^Qu��{�Bmb�S{�/����O�&u��R�3s2�E���|k�sk\z޶g�Eav¤�����z[o��N�-�����Bo��y[f�N�L�/N�w�L�1}��;1l����r9�&u �Z������-�NN�C ��r�o�t�s��ح{�~`@�磫���:gKҿ�H�9۽=��i땧-��Ё��WZ?��j��9H�֬�������Y/M
�1>Np97a�^�IZ#�܂��)1��]߅\g<*�NF�i���ѥ���i���		��~2�D�)�|��O#�٥���g_p�!�{�?
xH�*mq���X	���ܯ��ٮ9$��f2vh<�B�x"o�&N�|����]H���Mτ"g�ھY��{t\�j��+݄���^۾{8lz�Ţ�����6���\ֈz��r`橰ߛ��a4���x3���w��f������|7��_x��Hm�Pj5LE�)3֣��bF��buQ���"��jI�t��a��jZ4$�_��L� �&��)@!��V���� jG���D��\W8�I�H�'O��J��P�k��Y��5&EJ5O}��XP>����4����GX�7�4�o3(=�<����&�ʽ��:�P�4/��`l�M�Ai����5��zϿB)�N�yWRKE�2��D���UA����!^�
��,�IL�U�L���AA�))>�:��O ͽj��������'EM��K��y\��z`i�]���jvB��I�H2���h)b���cU6�fI.:|���H�Qfǲ�ᗱ_P\`ɡ�q���J���%�#Ѻ��T�EZ38�����m���В�fu�4Y��;K��U�����<�A�V`5+�Z�Tq�g���-�0����|�3�%��sdddl�	�}��������2�H��� �/�DZ@�RH�_{j+84�vT'h�g�U�{�.��L���"|��O%b��R��x8$>�%��dUN���� _�y�4��i׉^����jk	K#���G���D����x�'����S�QP�G�zoTA>�S����W����Da�96>>�B�38c��J��P	
}��=9<
�P�E@΍�vƢ�w��	����D..[�T6��ZF��M�>Ԛ��30��/y���͸w����|�N�X�?��D���S�)���tݔT�t~�q�,P�_^M�d�q����p��Ɛ7�J�l�J�1�Fl΃���Q�Z�}sV��/��&���;�� ��V�C����A���֛LD�ԏZ^��`�v5�j�A��0��,���J=��>�I|^�]׿�49i #�yA��c�К�!���ԛ���mek29!��FWW��n-������d{�^C�
�M��d��d�L��C����]�[�3!@�������JPPP����D*����Y6�R�"�F-�O�p<�� ���ʽ�~������1��ߏ�@@A~��=�8��5��ɽH�w%�A���u�h�͝�s��8��Li+]گ��v\��Z:0���4t\9�e��y�;�!f"��n��Ҧ��M]co�΁�Qf�� IEe��^�%:���1���=v���P2�z���sR��,k�S���oi �7#�"5���yuS�����qk�h���l���b�2@Ĵ�/C=��͠�V�v%i�6�H�cه�Ͳ�� ��T|:I8��Ii�9�B^�ϲ W�����������#���1�s>����q�c���(�m�6��~����|�DlԈ��"��jw5f�ez/���;o�#K��ϊ�P��}<,''Ǆf��@�9���>8�6�儞�M�����9*﹗3�����������R��W��7�#���1���q`(�]��JB�_)�&�ƆtlJƒ�aLa�BC�\��$Zs#�s���9�ⵯ�3�Eޢq4Y�)�³6DTGe?`���p��ww+�����7Q�fЎ׻��1�9��%U%�1�ͰO����.$�Ќ�6n��~��37�9���t�w3�3�|���u�{��g���9�0����� ��i��>��i�D1DS�9n�!vc�:D|�gmm8���4�@�&Ad���dH��V���u�w�Avw�6���+	��*�Oϝv�ϞfV$�a�ӬT*;���w��3UD/0�Ư�
������-���a�������ׅ�i�O���g}B��G�DE�ϙ�t���u�)Ն���>���uKិ�	����ذ!�!���7�?M9��#����Ĭz��eк+���[��Zj�>f�\�9q>"�"|�`��UB��zOլ�#>�|�STDqh��������%��L
'ӛ�� /ݙQ`��������~?�*�Sd �]��KU�5�G���:�k�U�������?��!Z�a���Q��2/K�7����+(n��h!:�M��Ȱ�n����S:�_��Ϝ�'V������@����#�q��RQ���yО8�uC�NN�Di"O�K���O�:�q��ȟ��(����ơT���,����Դ�=]r�/(AHfFE<�����*3ȋ��t�<�la�;���XX��LL0x�������*���;!�}S�`v�@ Z v�U�q.����T?JL�]5|�d��c0,��PF��<#���� vX��w�\���=_�ؾ��ܒ5�ǳ;���v����"4��9@�	Qީ]��mJ_w��%�o�)�v���Dk� �DUB�	W����.ZY�0.������Ed����~ ����5Ʋ�e+�/V*�҅�>��2��Χ��v"u����8:x\����(@|u�����X��C:q����J;E�Ó�˱�]H��H�/��U�Ս<o�D���Y�t����t+��)Z{{;�W�do����ӞI2���7 ��כ���SnaM+h�wa{a��d+x`M�>M/��=`��|)�ʯ�1�%K����d�����g�b��ז
����]U�{PZ>?0-c|@.�M�%a\zVo���x�v��#��� �<�=�'�|�xUv����%�t)�[�Xֳ�~�'�I(����.h�64V+�XN�b̋zˈ�)���@!`��ŗA�x�:����`�;����贪���=�{���;vΒ�Z4�e���Lpp0drrr��<�N�{P ̎��zS�������Vq���PԿ�ݨ9B|���k��wg��3�TN�
z�-� ��7M[�+�����]��5f=60w�`�\6�B���K��y���	����w)%mIky���<j_ O��i�d�E��qU��@f��/��c��)����J����^$
���s��Zc����pq��Q��� �[�N�-|m
��x�$����<<vD_wE�nU�66��Ӕ($B��� #[)�뵬�VFCc��hZ��\��I�yV��>���b�Bs�ej����<9�P{|WP���B�͓�ǉq��9p9�5������\@O4��^�(�� <g k8�˧`�i���j'����)o?��(RM��f��$:����㛗��p�C�W]Ԯxk�G�n�����T���Zt�l���>�#]V_�hFae``>����kyz�{��v/���[��U��5���#�Ѣ�ȡwvv|�?](�����Ϳ���~gboo�ߛ�h���+_V^.�.b�����΋Ȅ)�0��|��X�~�p<-�Q���#پ�d�xr}E{P���H�ɱWH�6��Wi����'�$�Z�({#�/����!1�F���_���A�5��'>�!Htc'S�o�J8���H�)/���!�Tɸ	I���:�
z��ja��4����=};��aז�^~��V�ᗃ꒎�u�}���(L����Is4�D�&3\��%�����zZ���ӟ?�^�[���u��8�Pz�y<>2[4�8'd���c��`�a>]x{{{e��WG��!�9sF�}n�}ؕ1�Rh���BUW:"��X��A��d=�3k�� tLZ�${�8<�������F�E�)XhB&�'3�q��H�a�[�
M�k|y���54����z�������>�yv( %�؝cys���z�����C�����0N��sT��:���'��Y��*��GrYQ�_1��'Y���-h�R�����`���.j,$����I�U�lD/���M�!���L�'F��o��2B�u���T���j����5D�(ihH
HWNc��,�@�i=�tH�r'v�!�s�5�%�Y�f3Д���f��/>yj�&�8}���}��f���A�Ű�bئ蒨���K�sy�pB�3:���?�c�9]B�S ɝW6Dյ�:�G8��U�k��B#��>k`D������r't3x���c�������9��.�G~�Z͙����ɟ��^0��l��?B7\����/Y����s/�Ϋ���yd����:�.��10��Zn��ۓ8���F�3���|Dݟʍ�����S�u���p`;إzީV������	�Ԝ��w*�t��:*M�ƀ0�>��#�+��-@n�ED)�郵��v�9gU=ږD]y	�]Hl����g2�N��N,�QB���E��;�]��=���dȃ�,񙲑���Rj.PpF��5cr_N�����r|�����׶	�b�ֿ��٧��!/�^�Y��n���â>T�`pbbb�n>Eh����ˡ��(�O	�i�='�?Q`��D�2��ǑE��ڧT'7Pҫ&�h@�/0�PZk�<)�ӎ#7Ð��s�b�(���&"���� �6��'3�~_���U�,��h�f�!����8o��`!墁Y��H���X�Gd3o�eA�Tpq\���f=�j"�j	���4B�����{8nr1�4�.�����#��V<��s�9]����O_w�v�](�S�[���\����P�x��f��w�VW ���� Vw��}�^a����DJRF�n�*�0Bz'p���s��}�{#���)W���S���>p(�����;�k�%�<���q�œ�kz�!�^�8j��6L��*�����Q�W힮��<�R忷�K�Ka���^>����G4��lAϝ��FC�S�� MDFA�sh ��?�ぁc�l�����]g�$�����'���M���\�:� �1��������$��O/º׺�[H�]U��q�5�W��V�؋�,�tO9ִ�c28��m~2Q�"hHl���D��r��	/��Ps�[6E�c�����f�~��@�5i�u~{�7;���s�o�w�A���v�Ǎ��3n���Y7�>��MM�fQbCet���K�1EB ;��([}ٞQ��<��턉���)))��J�0�<۽��3�I~~yYs�.2��*f��_m);t�etl;D뉮�U�r�^�ȺsV׃�I�M{�`��0�k�t��ž7�'@�߯�ds�y�T$FR��*J¿�L$����E��%�B�N�1��_��?���=9������R�ԑ|�b������ѐ�D5��M��nGjU������������u��T1[B�eڟz�LDQ�ז��z��]ҡ�1�Ϋ�x�tʞ��_�����ڙ��]�v	�V�P|)N�H��<��p��#q|�d��2����t�gl}f*�j��X��������gE�%��Feuu�a�0q��W �aX��Qs�>c�f��p��:(7��-�w��59����JIO�a�"��^B����y55�>| ����S�?�ճ�V��Ċ�z�\��/�b�T?!�rN^E�H�Տ�a:I� �i�40�@~�Xŕ�d���Q�hs$�vb��Řl�e����)�w�y�Vg����K+�HZZ�K��j���3�X�SѨ���1��j<�(�u��2��� `������<����4�#FM��)h�T�x�g<�����!���)�F��!��z��Ly��QU%+M���,py�o��,3mS8��I��JU�?=�4	�8��"zLZB��W�:x�������q����^����i������)G����g�I�55!A�5�8�%S�+*T4���p�u
��-�UPPf�b��E�:<��(��jf�$�/���a��&�Kq3�����^��Z���6������� �u3�7���"����$lmTg{�OG���e��Z�y2�y�_��Q�q�qwx��$JB����n�+8�xՍb)�}�gT�F��k�>:w����Z���������w��ON�>�!�k����%�A4�=�����Ynn���~"df����(�#���؍Fa$o&V�3�	F�َ[��9���!:
��yo��y��0���|g�3���u�*�N�a��>Ƽ9/k����sS������3�ǁ�F���Q<h�.�=�nOX����y���;�'�{�	�u�]D�K�\$
�e�K��Z�*�z��j7! 5l�n2��ď��^;>�i���21_� �j�^ ��VS:7A^��r�3�7%�?}[�F8\Yʺ�TK��;f����a���%��5X�C)��{��_p���)�HG`��S�ۖ3�sE��[�䷴I��������Xtn���"�s<�҆��(��|=Q�!X�ń��q�l�����5C��tn�b,ŞE�=:�]��:2e�Qlh$�'?~^�-O�CeK}E9l�z2�~<�j�z#�jopF4fcbddd�^�J�_@>>���=*?Ñ��tzG�ab`�:;C�
$�2Q��4B??�o3��`�����4��E/8Y;ڠx~Qp�~{�#][�s��-v �Ƙ0F&��6;&k�b`L# �||�F���U�t#Q����ǧw��:{�y���-KjXtʂm�liv|�c�P��&��Ev��	��&N�ay�o8��*n`��.��#5ޠHxpn�I{���`L�Cx�����8��@�/v�Ah<��i
F��\�|,`��S~:l�T��%Pr�*&�:P�2����ôQ���j����[R�	$%���$͓+Nc\I_n��me���xC"��w��)����,���h�Ca����QW���8bU0jfY?�!:D��������=������9E:ં�H=5U�R3�>�����`�ʼ�N=�dO(ñ	��q �RkW9.�4]������r�����f�����e@W՚հ�i&�nEݣ����{��ڌ�2읙��������^v�)�9��n��y�h��Q_�-(��fT�5�Iho#0��x�'�n�إʦD��L�:�Xr��GHt��c�U����Z>V�~�ན�<�]E�K�r��pi����
e$�4đ^��K���js���>*�Wڕ�B���w�
��I8o��)0*���1�t�eX��2�$���/4�t)�K�_q߃5sJ>���.���������jXW�?�>�D�ؠ3t�(�"��uC,!r맰��
���UH��,F�g��\�R �Bk?}�ܓ����|�N�������_��T��o�5ۢ�(5�'"�t��U�[if�^B-|O��~�?�ǊzW��AtX�j��:��:��-������8��׵" j�(���Y?��鯇�,H�g��� -�����˞�j��Q�^M������P9����:��3��vG��
��*��r�ݦ�z�D��;V�.�ipl�R�zD��΅�7�tD�w!GH,p�eT��/v@}ϸ�O�nk�L�&��?�k�S?7�}<Ԩ�Y�XdN����l��-:�����<̾�"��G��%t�;r�̇�fp�V�oK*�b�;.�7��Rih�Ǧy*����_j-�U�@,��H5K4h�3&�!V����P�ˀ��^��"C�Jo6xć����y��Ҿ�~2mr��s�^��r?0OR�-�ܤ��;��9b���Ft�$�\��F��@L���J�M�JC?A��q/�7�7���6�ժ˥j�ء������*����M���	��_9-�P���-/j��v��Ư�����Z���<s�kD(�@��p�:}�5�sE5���\"z�V�B��éu~�Y1dTIj���Nv�v}�f�</�nO'8H��.�g�}�S�6_�L�Q�I���c��O��;��=�:k��Hd���x�yu7��;LKe���@�TӍ�۲2�`�4AZ����~�,�;=��Ǹ�����%�	�x:BZ[�.�Yp�Y�#c'[�L�/AJ��H�g!%{�޴���x���	�ZF��������ŧ�2~	|ݗ;�Wq���'����&���)�=��&숃˺���r�������kד�����N�;�<�]&]��kؕ�������j0Mf�Ө����o�+��_7"�6ɪ��>PxN)����z���=�W�r��<�:�:�N,-��l�V����.a����ŇCR֭]�Z�v+�2P<�SGYƕT�����d	�#�;<s��nu��/��(i,TA��P_	��y�jV�`9(�9w�|nC��7�깂:<�y�����F_zot����(�s�a�4iJ9�{�C���fe����G���;��W �=s��o��pD��{q7��oGz��>\Xv�zY���i6#��6�}M��7C=�X�z�i�}	�L��C�,�.R�@��I�"~Ґٰ�s��mU����:zh�������Y�Ы�Ԟa��fD��$��r����}�*�~SQ�Ϊ#� ����9�(w��GU�F�L���9��'N�f������߽�����[�ڝ5�CPX;`N5�b�㢻u�ek� �*��;��%�����j+��z�k  �����/M�a6���U84.��g��/�{=�	|�6yF#w��2z\�ş~�T��R'��I���Pz"�AH$�1�H��/�8,ںF( �����E�O�)�^�6�U�	�;��k(_�M�3$J|e���d�[NVd�-|]k����u5Q����s�)���P��;uD��Uj��5��v?���n����ا��[�RS�7|A	��1k{Cd�ޓD���s*4L|خ��q�؍2�cC�V�y:��6��+����k>�b�G��)�hh$(��WC/�����Y{�,���)ښ�q��t@Xkf:�i�P]{��o{�*:�|@�?��>��:h�*�v��l�h����cGZ��տ 3�'�,���F�Q�ۼ�����x^�p���nE�8���c�`m���Y������X��C{�ř����[�&��T�����틳X#�O"��%3��+*X�㵩�ڿoۏ~����5b�`D�U�������<:���[�x�^�{R��.�����ѹ; p�o��5�����WO�����Yv1f�_��,Hx���V�f��������x�tL���2-lX>x�W\�^�M$\1���>&��J�L_l��&�f�'1$������=�P��0��~)]a$.c}(����ȻmV.o������v��#J�!����:��M�o�o���||	f5n�B7%����i��}Y������iv�MD�7�O�V,�Q�4��mڢ���@6��wֈ$D��&Sjm���1������`9�S��l���1�g�'���4�$� ���wK�y[C�~�o�`[دܱ�~�?��D��y���j*vԜ�e�t��8'��s���J5~��޲=v\���~uI�K֊�O]@����u���G��$;�x���_�!Z{B|�������TPK�$����΃�y��d�i�:��R�O�xlwzL��S���~b8��]5���2P5��b|���Y��lX�ST_K>A�Ɂ�+�
]��f�
��FdK`u��|
f��hg�B����l���E^_7�[�\��xz�H���:���^j4��k���s�g~f`N��Z�^���´��r�G��JU뾢��D:S��;{�4�]�B� �3���p�[Y��&�j۔Q����O�VyT�yt�e�x�x�jl�3F��{������ߥ�s5ǟs��	���P{�ޢE�c��9Mf��z����f���/�[+p��A��Szaw?��A�pa���n�ƶ>���i�V\����o'�k�E�W�&��e����)N(�d�Q�rL�Gk_5s�iI�=}�載`�`�E,�N�%��]tw��矶��Z��_&8���<g��[^@5�I���O~�t�6O��찶�\��=}���7����uq��o߷t�B5�z% 8?_Rk�}��)�c�ZG�1�����`=̇G�\�=6-����"�?���[��ݗ�h'�/�M�_B�h�N_�����A���Uu�T����"
y[Ջv�iI�w�b��g�堙���g>Oo��kM>ʇ(t�����t9^�"�k�52�o�y��?`
�?�q��K�)��S������.&<��0]�KB��L�Q�ve�Y�����ԸC(5�g��Y-fTpN�@79������xg؉��%V������6�=���h)XǢ�=��*P�}�ir}�$b� ��e�\�3a�ץoG�/�R���/�'=����9��ɓ1l��N�X���7SO]��j�p�6�j%����2�T��W�?��G����I������bF�nzH�';�!Lh�i��:m{�D��M�,my=!*y��x"�v�/�:T���,�;����4���YҞ���p6�mo���o�z��[+��˱�&n^����M;���/$0��B�b�C'[}�.��Q�2���πS��j#oB8���N��~�S�p��xǒ"K�p�M����XjD�����6̑[{�Q,����M�����<3�\���@|����������N��*\�(������R��gC(�J�3�d9�T�~�U2�l��/D�?�5w �GS��{x���69��۲Vdol��d�qS��P��RCX����HW�o8�7�=*	����W�>���b$*wpr�}_u���QE2-�Y�z*f���8V�Q�&�f?���OǗ���d��4�Dsz�%Ζ}�Af�_/�#�S����R=���+���F&��1fx�YДe��tF�FĂ�/����:�ܤ�@=υh�FF��=μ��6O�r��}�Z<D8�S���5'Th�3-��	�tǾ@�d����LpWD��ՙ	��)k�H1�	m{��cWr�u_{���N<��+6�l��xw�[g%Y�k.�VR��V��&|�<d�Ώ�U������D-*1�<�,#�7�t4�y0�a���ʲN|u�lI5��lL��~����ͭO]	���S��>��V��=E��m�Z��}68Ǭ6L�}�����a-_$F�3��W�Z�g� ����+-�T�$R&xH~_�$�@h�!iQ�e�Z6v3GJ'좊���WҢ��m���{����-ܠ����{�*��Yˮ�:�)����Ӊ�?��K���芡��ۭ�,����� zy.�@� ��Gs�+C�b����[�hf�x=qZ��^]�'�/�$����}Z�_b=
�I�ژ,}{>`���TT�cnКɃʿ�|n������L�R'�P{��o�]_+Z�AQ��7�ny��s���t�Ã;���!�wwwww����݃�&�������'�+����a�T�޽W����>5��b7���Z?g�켯>m}�$;l��G��qo�O4;�E#>��r[>��w_�h��b"�Q�C [��[ٻQ�D��⯖W%��u�n�h��	�O���G���D�Y��R{ �,~p��۲���z�Ğ�W,]��=w}����{�f�W�]Ix��6���U[��5���gN�!6=���D���\��� ��O�I�@ű6y #��n������60P>�wt�F	�!�j裂(�P��;�D���ި�������\Kџn��,��u.]�q�f=���=7�fQ8@D��A#������t�}rq�U"�	��1�/��a7����l'�3�_�ZGn{y؟?H�}o���u���@�/B$<�r�m$��½���Ih%ڳq����%�ɢK�43�m�y ��+����m�v�/��X�Kc LS�=���hIG>Ǹ �j���>�Vs�����-[�SJ}4f���w��ݬ�00�&����ȑcH8}���B���&M�����&D�9q� �~�Ȣo*j�Y��df׷�K������zv�:��]יh��!�z%���)��v������p4��<.��YD@E�(}j��y�ג3��s� ��d0]�q��BF�tq�XSe�s���1a��J~c�'�]l}�=�jh�(�n��j� ��c ����$���,Z> r�Y����m�?�l��3���$ad�;�aQ�w *�e�>��Z�� ��~R���1|dr�}�)onx�?��^��Ȼ�T}߽��+]���'Տ۱�b��s����!���m��(���pZ�u�e�H�9�W[�F�P�������JB���N�3����7"�I��6Cn4y��n�G�8�|�y��|q�a�.�y˸'^��Ԏ��{��о�VB�M�hb�`��}2�6SU�u�1 l4��h��%�{�>���2m�Hc�l��F����F9+���̲����d 	~�̫�3�"ȝ08/�Z	���ʱ��W�OZ!.W������W�Y��I�f���H���@A��T��#iz�k�t$�����eVPh�y��\ �%l��h$����?V����	�j�B%4���z>�U2�M��9��XI��i��m\�x�:����Ā0��m�hv����⺦��O� �]&��~=Y��f7��X,�:s(��&�i���؜��#��:��"�*ǫ�OK�>�O�͸����ZI���>J�݂@5�x�6��J�^J�\�K"�1�e�M�
c0_�j3�^����V_�D�	S�7J�1R��ń�]&D�q��ڥ��jrw,��t��|�r�������sPҎ,(�u&�	�c�DM�j{Q`���wt��a]i����j��[Eؕ��+QVÎ�Lr$U�~Qm$΁�V��U %"3#��o��Q$.�Ly��bƠ$@��2��l(!��a���;�c;fN���}��'��LN�ciwÁ�������@G��~�jO�7ƚʬ��P�>.�_�r�j؈yz5,�͟Vw����$�{�T����Yߖ���,#"�l��m��2��o!.�ӌ��G��,rOW�2+�P���jԦ#�V:��j�zЮ�R��}��&�(k���k���\�s����5��'_i��Y7�mI�R\/9�F��>V���>�P̿����x5��	0�	(�{w�$	��Go=��*O�y��>j$	`9�"M��̼p��D�ˋ Q�Or��QR&���3�â~�p�d�V� 0:�Bo�[�h
>4{$@'�F����|:�>:V8K��{n�׆:g>qz�By`�>�^a٧+�q]����[�G�GM�IR}��G]8Tl�����ߤh(�Q���U�"a�1�F���PB�p�e:+q�j؅J�����Ћ++G�
Nf�Y�5*�3<&��p_tɍ���U�*��mMvS��k�>��I��u}p�
n�Vt���Aa���]&Lц�GC�:%d�Y��;��˷�������{w�z�
��O\ywJ�o��3f�������#���#���pj�Kt>��f��\�P�X�L���zҥj���YY��1�,��L�4f�cG�͞��!�7#�m���& �`?)�!ڜ�1?v[�,�Y�Z�
�<�ƴ�y�:t�7��/8k���M���p���**(��CF/�q}���O�)ID�M/���Ǜs��A�&���Jo#$�]��($	��ݻY9��$���n դ�IE�sC�O��q��q糶�49������� ���9�?0���x���������z�N� C�Y�p�����I��~{wYY���r̰qд�-�K���F�ۥ����ok�߸�n���ͬE��k� b܇�%!��OIR�ifb�]� M��F��c�
�T�fs�$@�iXM��7T<>Hy�2�d"B�.T�~���;�:[:�������3��$���H�Vpp�]H���=%wOFR 0ٰ�
�u�yv7��j�#J��Ng��I�st�륈De��ԝ�L��X$5���������� 9 \�X�
�Y��0���})�++D��/l��֪&̡L�Ύ����7� �cD	;m�ޖ	w]��)��%׍b׹ݣׇk��
�\��e�� �@�Rw#33Jq��Y6vv��Y.;Εxq
J�Z@A�p>�|��g��"C
���#@�<<��-2@�k��y��{�NdEx������=2[��>�"���U���\�;g=��^9p�.Vn^v|��U�*��v̅��SU�)E�$.j��g,Dl_�|������(Oxb?fL/�s.�����jI��=�����S����9v��1�~C I��uWǷ�g�ӎxZ�����fe %�����`Aj�s@��8���&��#�ƪ�pnC���tQۀ@b@�'hȓz����_�Rc�����\��6��~�C��6�7jY����\�0Km��^���o�FG�'@`��~E>2�U������n����?�;�f%,l���OU����_����T��~2����'�AG���Kf+ʣ�ҋ܆�cS�����I��%����j�f���������1]4d�N��+q
����&n0�ҙϹ|sӃ�̹�tQ��V��W��>6\���zCy7?2�rn V��?B�ў���aь��E&͗q��]ӫ:�@��5?	�I�L���>r���\se����q����@E(�`Xf�J" yQ��j $u�}_�t����QϏ���ŝ*}X�H��e������&z�eii|2ev+`zj�ב6���j�+�έ��vB�iw�&��s�ᣀ�H����'�q��Y�A��}�YXu�Q�v�;A�x�Y�����1�f�+\ ���	;,ܞ#��+�˶�}����6�
1�t��Z����M%�d�ڷ1:���2�2�X�W�#k �UO�rjk�*.�fJO�
Ñ7W"� ]�0�k-�= P�?� � �O�=��O���cwY��6��̗���R��V�Kx�h�[=5�Ѽ ���>�d_�+�Y����Mӄ~sC����<�:MیnÅ�$��';U�����y#6$]t�8��4kP�R-j��g����PWCS�����;�����l�<V��vsJ���b�G�)��h
?����MU�)r��P~92(7��xbOԓ�7���(0��2H�|$�Җ�i~�����^!e����	566����O�~fH)P��O������V��6�����@�f����Q]�ME�ܑ��η��L�A�<�Rp�Rm�Q�@�
LQW=I�T��|��y�n�����yk)v�i.&�s 󱷋���:�������tA3��8�>!*�Ĩf��p[�J��N�Ξ�͞6���t�3e��#ƚ�T�I��m�ًf�v~��C���w=���Ҧ��ug�C-)݄Hv?SN:_�-�s�Ud����~O��ܞPp��z]�(v��Ŗ��ǳ�s*��<��5����4iVm�5���'�����C@t�JA�Ƿ�-����NK�7׭���Y���eS,�@����}��$3@�p�_Y�>����5�����5ɢ)L��\�d��3ڣ��� ��ᷴ;���0 r���,te�N�8�}?���5�0�5�2��} �=J��y=�y�b��vM놻ǡ*e��#����M���J�40�	�9�4�žzt�A(��!���={t'�qfw��{��M�
�-��_m#D<?�1��MpTE��44�~�`�R^p��I�w�\dB~ȝ=�Wý^���c���!��+�VQ&���bv�1�����#b�,^����t?�ǆ�&�a���K�WE&&h�l5����U  ���q 9U_�M�`
�ؚӑ��'�]L�'aU��f��\�����*�'�2\`^`$�w��>:E4u:��-�L$�F�--S�6���z��~���!�A��=����)xʴn�ɕz�����0P��I��~��˥\�n�K�4���`� ��k��e"z���{���'��͆zW�A�]�N��U%�O�2�Z�Q��(b8���In17{�1�G���_ T�yB�8o�L��s�g�!m�B�����Hq�E�T�_Ru��t{!o^����ե�G)Ä����BA]+A�Ct�M2pE#FX����(~�˴���s�bQ�-���׀� �
�����?280[;�c�G������
�h(��p��D�o��2���U��T���T��)�e�P��\iݹ�S�`����QN�"�Ӕ� y�ڇq��җ��ZDT� �'���őۏ'��� �'�L��^XȄ��cFQJ���5s����R=����	-��~@]56��.���bd&��(fE���Y�@��F�@ ���UƯ�#�.j@��
&4���w�߽c;��˓��'-c�w�a`BDb,:a�?�3���y�W������+�*�'EJA�6dEQVW�a�Y�(�aN��j��*�~d2�t�h�R*ּFV�W~q~�HOvx�I7��'v��i�0I��`�U��A��7ɿKY ��q��~'2E ���;�EM{3��������&{�.sƮ�e(��@xT��@�C������;��4���SI%WP���F]zZ�5L�_k+z��N%~�3A��[�8�{M܂�x�k �¯2RpJ���X}���XW�d���e|+�W�����_w�I���/�=B����˩�C�\�*���ږ���by3�œz 1l�@�4�@%2Z�a{�|�gU�}]�ݷ��$D�2DD�;,�D&E%�^m��wD:��u��m�����&U� �'K7�����23�z}5�h�(���^)]��[��'`����{����m����9a�j�՞�����/���/��u��-ϖ�lQ`��|���8��9�x��BL�P�4�.�x� ކQF�JN�5�U�<%죙U����]�"�� iN��C�5�n�u,ځ����.eD�˩���y�F[����OV���TM˄ԎO��]�7{k��T������Z��I�4{�!]�7�k[s�M��0Nd��/|>�k�G��1Fs�Q{�&\	'�
����T���&�_����:y���:�9���n[��t���5J��a��dS�XǼzA��{��Q���!!_��?����U/�����!���ҵ�U��Ϯ�LmQ�ĝ港�/�T�ZoX3�h���M�
�(��V5g*�iw+��Ř$G����P��F���`t>�`��;����A�奄�����t�x5</Κ��KX�z���F;|9+���*���f��	k�e��W�2�Y�ʺ>�Q��x��.+ף�)
D���Sz�����fP]�=O���ּ�;��1-�;^/t����W��<�w�=`"J�4��r������!BMA��B���������J�$w�	�?�iW|��a�kj�x�j�EX����9>�������7�i^G3��i]�0Epeg�q��V���p���փ��%/�:[eg�<��;�o�7�1�E����_e1n/��5S�V���*1���ԛJϹSB_<喚2�S�"��>�!؂8�9U:Ci(~DEZ��V���k����W�,q�R$��u����62t?����Y,�����]ɐ�e��u1UW0�m4�QR��������k満�/R���	�}H�H�������߀�i��Q�d�0��F�"
�L��a'b1 ߸�|�C�I76Ҳ��N\\շh 0����qft��O�~�VOar��Qj((xtt�Y�=���H�Ï(���0Y�D##�9?:��!�w��������kr�Y��
�������HD����u���p������~XcM��ˆ�]Ƣ��5��k����v"��5uT{��Q��_4č��:CŁ�I^\3��b�UA\�W���0f_M>y�_�c���?�~�byRc���Z���_�m0 ��c�hR�~f-w_[���m�βC ���f����w��z����Dx�4��9�¾j�,�h���a��`���pH(��"8i��A"ZW�*��&7��|��Q�D����L�23o�D��M��D=�xFˎ`��N��Hw��8��<�B*�olɔ�PT�l��Zs/�0�-�-�}�+6�-17�ˁ� O5	H1��B޸�!Vm�+�]B_Íᱟ[����o�Y�5��o<@�X��}@s?r�ˢZ[3L�#y�hzV6��.�`�c�NY�#)Vp?y�豂΍L�K��8%:��S�\H�l^IЖ�(��Iu�6�f����5�`d�JY=��P?-��Y�ym\��R���+\�O|����x�x���"����p������o3la"P�����/TQƽHIΣd�W�ح�Ș�1U���Cd�e��� ���`�.x�B�U_�b�9��Z{����y��z�z�.�d����Y��@�?G
���u|�VO�CUGЦ$�*Y���}{m�����[�ǂ�;�5$Hm��ڢ d�}�>D1�,`6���3� ��(? ,�h�hvˢ���F�e]�aH�\�������|�,���
maaS��<y�IU.��������0v5_���ݧ�d	q�9v$R|drqӒ�x:A�� Y���1��(u�R���.S�:��Ҿ���4W�Y���Cl�EVF
�U��^�,;�a�����"e���~r�D�X�E�0x��1Fb��xvA�	�֭�&�R�Cʫ�I��ԏ��C���h(J�<4?�O���,�t�90	�,�3n�SVY	�f�����v� ��͏+)��DB��:�0x�s����хQ1t+�V�YVl.�4fO������RQe/�w@��2��@�ؠg���s�s��|Q��y�PɊ�w^9:�ve��´�2z��2����y�߁���9l�0�K؞��
˜�,���ۈRW6���:R!Rd�qqj��IX1x�ߧL��PN8#o��AV3����4#+}��`�iW������ks��z��L�f��PR�A�6���a��zl�1iۡ�[9NଔQ�?�
6�0cL���y+��I�jd<=xTgt�	�XS)�����nI�Ľͻ���(�P�X��DF&�?���b&A\=���S����}��4��s6ZA@Cq�����S��~�ȧ����}�y匑�"K���䁫�P�Y+�%y��gsU�,y��'W���	^���+]�A�s+�(;@h[��5�]��-����[.����
����t5��a(CL�^'��	kL-�u��$h��#��j��g���:{�p��h��?�ׅ��P����kIL#M1�Ч���g��[MG�f�:���3�����]���6�<��E2
v�R@�;�N�4��~�WM9��PK�qG$�u���0@�`3Y.%7����zt�yd���-'n����4bO��A�Gԝ���*pG]�tD�a
P8:�@����ɤ�mg��@)U��	�^�ՉJ.җb3ԟp���5����[q�6G.�6�&����ܔ���Mn��������M�dV�y/�E�b�/t9�$W��Fz� �+�=�I��v����H/����94�TC�}���i������{��G���6�{`�|��W�	헠����!/"i�c�>�*Z*�w�%Vk�
q���d�L��{p�n��`Q�C���4��dɠ�Q#�{�s]0YA�7�)!na���«>r��bG�KX�.E�~�1�+ �O����͟j��=&�j�9W��D�|7��Ф(�����s/t�
NA�9�S���)��>�[�lu��o���ڍ�bo�wV�?o�/�{�U�����z�.��>̮{���5E��n���"7Ҧ��r�#�#Kj���韖���P��u�˥�H�v/_���uh����m���t�`hP)�#�]4�z����{<�����8���V�}�����p��4��c)5���HfQ+r(!�J��</��O��?��_��;��
퐌��w��J����i��.��H�X.z�<���U͆���y�����6	��m�K��.��NGc�%=��u������ �t�%7A��ZÍ{6�Q
z6N�`����@�J �E}�L���jӛ���,�㬛if�I�T��Z]tb���v���×��ڶM��9����=��{2$�����
)��|L	�_x�8�ѷ[9k���Ev�M2�h
��-�5����Z��KpyE���t��C�c]��}��� �A��/�>\�����C*S�ʯ����)�;p�~m�A8u桝�6£��W�Ȳ������T�t);z�,+��O���������SC���iנ��JE�l�Q��9޶8��{�wͯ~]tf[�e���f	1�^�)�z��'�Vm�
=@^��g�P��6���^��c�:v���kt�~$7�(yE!�$�4& ������K��(����ӳ1wo�C�}�j�'����!F��6s'/���FًJ����_��	��#���7�E| p���kpr�ә�!<��I�������8��R�v�b/��N��p��	g��9ݔ��BW��B�-��jQUɡ^K���ij��#��ֳ�掠�i�P'��?MmE�ɬz.H���{
&M!V�Ԁ�
�ޤJ1�Ox��y]윪��o܃*�q~hu���G���h�_��s2��I(G�~]p���l95g�ѷ~�f�Ao���d�}�����t��Ty�d=i'��
D�����~�Ot���m�5�3C�0~�Ӡ	����E_��q���������J(@X���C��Q��������э�RL�{�pR�?�m����z�	F�l�<g��Y�:b��z�,��z��ϟIٻ����W�l
RfC'N��n��l�O�|q=���9�'�_(���x�E�^��=�}����)M�&�>��V����pc�}$����]�,k�O�f	��PHEz^��k�%|*����	ȗ>=:��4y��9m3$��+P�tH��0��F73ڕvB��r�nZ�Z�?A�R�۞��~-ׇ�����hQ���/D���F������c �4����A���a��*"m����,���r��3~K��t��IZ�.�^�5�d�r�y�U<�cx�-!�����³���/��ll���[�;ރ+�����/���h������/��+S��u��8���|��vNS�����e�K\	^��]Dq+�m�A-�3�1�8��H�hd�����'�cRIW��w��&�������Kb?�^M�5mO_�?Ś��'������I۪�������<��惋�J�
����^�J�q�[�Ŵr��B��[al�r��Wv���ۧ(sי)��?~��M�#�U��ik�*W��_^+U� b�F�#`�n�s,Oy�ӽ�����r�K�"ZAʼ��9(z��� �!}TQһ�K��n��E��e�@�y:W�������~��{v����n�����Xyϻ�3�� f�.�um'��ٿw�����7���Q���UZ��߰�������b���c�#qt�
�~�&�u�&�4b%���u}ǣ��:��s4���Q���ٮ� �1y�+�s���[�<��Y�Y)�Zc����*�᠙��� �:z��N�;��Ңc��ID��Ƿ��7Iy܎h�7�~�7GT�B�q��D����z|)��<_��O~{|٘�!e޽��KB��9�*�_�'���.�|�d�NԺe��0Ns51���S׹���ϫar��
�T��h
��h�l�i���y��4q�8w
^6��o+#����w����V}Z�	k���v���Z4m#���+=e�������̪#�#���/��|}ص�4�x<�G��
T$|f�s�z�2M	���t�����%�����Qҧ�A���MQmJ֣E~jаF,�;��nq?H��K�f��#k���.��E�G�p��ǿS̢�}��4�=�%��9�'�sEm7&�n�MP)���M�nF��p )/�(~h�k��*����FP�-h��B^D�!��ɧ�k���� e���l�A٩�7B���a�N��_�Ub�f��l� ��Oo�\��v>*��h��.��>?"�܄�b��y[�p�����Q|�(_��7����3�=�?�iy��zo`�i�Ik��:1��h���Db��G���8�_��nΐ%���q���������p����:� S����L�ó��$�?����hkϻ�x�󬭷KG /���U�M�L��q�8j��EHv������k%��X�>N��@[L�fRB�J�K"8��qM�*Mx�����mܫ1i�a#�i���[T҃��;z�o��j!)K���1��f��;���U��t�>	�Ed!�i�U�����VR���aV�$2�@8��+}#]u�-]n�����Y��!O�G�)o�����v���p���&o��[�a?ҭ�q�1����9���N�5ѵ��C��6�Y>`��~-�[Qn En�O�[&��I�!���*���&f��?k";��Os�Wr�x�/���DL��7uC�!�2�yLa���pNU���E0ϛ��T�޿�*��>��-x�`\�}������qN�x��	,��ߧ=	�L�E��u�p��-^t�Mw��f����ز�]���_G����"�E�C�Δ��7Oã��+�J��?�[�K�Y�4���xp��ٗ��[a���R#��xB�/R����I�/���L�Oa���&~ ��j Y��C_�HH��N����2b�$�oV �*3��s`�Ê�C�UW�7,�x�=��!���?���jzlx��L*ZK
�+��bv.GZ�-F��Qg�e	�oƧ+��+[b#�(�C}H���6K�)*'�gb4���CA��q�\%Pj��TE�ol�����D��(�����h������i��� �m����14QV��Ens�����à�v|ﮠ�����G1�����+�������}u5��K���ٛ��n�����&�ؓ�odu�&��2�H��%��� �!�p�.:kѰ�ܨY%�u{�3��̰e1Itl��3��k?��MTa0���. Z�n����U���p�T�=����W
Z>
�	�#�o����;-8��=��&D�(O����V�� ���ϡ��E�I$��1���CEIt�z� a�r���H�F��5br��.����Q?���
�Ec��:�<�"R�zC5Um�p�Cd-��o
��7;��k9~����6�����փ�]��r�C�`\ �'����`t%ߟXV�kUU'^-u�ΝOi�n��Yx����\DT
�dn�U�,�X��]s�FN��$��!`�;�q-➛s����_�w���mMF��տ~R�ߠ �ˊi,$��U�N����K��B�c>]  �V��E�E#�l����_��i�&�΅�8�!06��Qt������>����M��C9-�ZY2����6]��m �*������bh����,��>'�Oz���z�$�'�"��ʣͰ�:�T�r	%8�Z���ZS�W9t}��LU�k>[s��{���|Sl?7���6�xH���cS�/���6�!����<�@����©z4.�K�����"/M�.Eᵪ����L�f�V��1����$t���rr���s���1y��'�dG�Wܿ�3�ض��b�A�jn�Y
kZ�df��p�5�6���;�fɋ�>��u�x3!��d7���)uրן�kg*�����(贵�v_�p�`�s/mg�z/�WUG�[�h4�MPh�D܀�{P�7!_��O��^�?O�W'ְD�wa��u���rvy(���y���HpbV4����ן&?G߬�a�@�&e�`�W�IG�1�u)��1��,�S
�^��`+^��%i�St�<ɸ`Pe\��|Q��7p��d hj�wi?��i��@(���y�0����g�x�5�\��V12�_�Fl,svw���D�_	�s�T�"�����7%�T�VS��v�U1�e���ϝ�Z��5+�Q�01����Z�8�H��BV�I��^��M��?�K�;��Nψ� �y���6�F����p��ʜ��-�\�
R�_��b��aퟣE��d%����q0H,~�p��K,���h�ݠ�(��A�o:N\`�8��W�Z��~����՝}�yk���(a	���@�_�7�	��g;���L՜�5es����E�6?��$S��`TwIS����GW<ϗR}ő ��L&��Y�T��4���Px}�� ��,�t�����#�o!ms``����հ�Ͳ���p�u��w�2��E��I��JL�Y��g�k����K8&����H� � ok/��,X�d���M:�(|�b׏z-�WЉ�Z;��!��T��p�DqHh���Y~c��>�r�<y��r���=�}�b?�qd�YJ�n�i�x4����U�6+T�B����_�6���/����r�#�Ut#>mWOӹg7☨6�=���"���3 ĕ����s�c�}I�N�PǞ�}��Gz�� w��1�r���H+�<�,�����kP%T|��g� ��}���bfj�{�D�$}�>�7?��=V�b:�g[�h���Y*�)@�=�exr*�څx0N�7t�j:��VH�; �│���m[�_xx��sN3b�t���$�K�Y��D���p�E[�G;zJ��@��ӌ��mZF�-�/�g�X�M��Dԯ߶���z�7?;j���N��}��as��p�^>,a8�-MX�ڲQ�,��S�:�O.U�<��p���̔\!p�C���wZg����AQ�n���Ǣ��."@��o�]�t)*�p�]ғe�.-i��?%�m����5`�!��i�F2xv{��%	��M���Aū�����3q*��e�|cl1��\��]��I�x��y�w��K��H��9�m���1�r�B��:���p!b�}-�"~b3e�����C C_
�g��/�~�i���$B�1� �M<}IsP5 � cb��7V8���׸~��g?<��^A���V�/B*��V��}�q�MyIc0À�<UD56��/-ͻF�y<��n ��HI���֙��o��z4�ᵢ�y�����)��O�p��������ǜ�����9bb�7�2���׮��!��v��J���5`�$�m��L��H��������������,Hxri�u}f1��Y����0v��z������J��9����)�%t��;�J�=w�&*�G�&���9�e���I�"�)z���y�M6�I���)�+�RI��]|QF-�rjB锗W�n�TL5_1�����9mUf`P�;=��  �D��E!�w����v����W���Cf�e"�æRV> M
���8���7 �w!���O��gFw(ߠ����5f�je �O���^�u~:ףj}����ĤR�.���4�U�s8oa�̀�zѡZ(�4�i(�_*
ܳBaAl��3�3������wP&
YV	9������M�D$0w�A5N�r}�f������zj�08QWr/D�+y�/J�����>�(	=.��puMC�d��F�=�W��v�(
�������Ks�$jj�%����bt��х�/�.Xq"��AT m�,�T6'n<|n��m��$`�S���==�ᆮJؠ݄�3ѹ��ܫ P�ֳ��BSK������<��κ{.�o�����g��O�yb;!QWt/d*T~ܽ>�8{>c���WD��h
�����&������*�����'���?pd�$�:T�\�g�YD�Z;ՕO�ȹw�k>L��&�}A9��L�	 B>:CǱ��� �
��C\�v�n��t�v5�d��OKW_x�����A5������5���YR�e�ʘ�=Y��C�|��9�d���`���Nm��Z�ݎN�H�I���C���ߋ����A�F7\/E�yB�O��p�̽e�"�٭/6	�
1{��\-�1*�w�^�ۚ���k3��]�)|U���Kڐ�G���u^�2CQar�c��?:�����X�`�՗�
������8�x�]Jl���:˜3�ޯ��]��ٽ/.�/��EWD�>O�<@Ά41��5����ݹ�-+W������.��'��>&��}V�,y�'��bDO
\L�C�D���2N�CC�� �����C%���H�X��C��7/���ߌy�ZN�͈�c3�����[����d�h��Pt��jD���>&��ϢYY]^@�}��2��"�Ί��)���O7{n�d�K�����Ј�D�B�q{A7���'�� ����s�$T�;���PR[��ş/�y�Er0�x[(MY@�"�"`��YF%6�+3L(4:*����J������o�������n���?��כk-�u�_�G�@�:r��K��F��z#A
)?,�I���&��.�t̐&U?��%��3f���1fCI��^��|���C�e2o��t8��Q�s�~���d�"NrA�8�M��䷲�T��@�ϟ�١ �M�?�H} �z �g`��)���5�H��Q�o\�o4���B ��fr}���p�޹D���@�;�:Kb5�tُ/���ۯ!؀P����G������b��.)�K�u|k�U]A�+��iv�b��h0P�L�@�|�61�'���f���R�|\h���]�BޑI�0�EԷ4�'ߞ6=��zPti|��rkF�N�����W!x��00Z�KX�x�|��N �F�#7��Bt�ܔ�<�U���U�E�_/~��mvz�Uiw����µ��XnnD�+w��f��������]]��鱬����"��j�q"����Z�hd�5��\�#�#��ƿ�q�+*��D���.>�W7��Ð�,�k�JNdu�3�S�*=���U�i��ߠ�q����2e�K����^c��f��c[�I�w��ã��њ�j5+�p�@�c��'���ȱ�hӑ	W�X�\p
:4DQQ[��F�J�A(ʴ㡫`�`�;h�f�UZ�Cg6.m�m�ͧ3>�ٱL��l����/W�;Wapi"N	�l]p<e�!�堖bwa�ݓ9'AA$`i�ﺦ���o�v�L����Aet����|��+���Ԟ�4yyEӡ�l��6�Ax�OJ,&�6�z����	26�3G�Y���NRB~�iv�z��u��}+)n�CݓaDMu�Q�~%ᢣ��D��%}���ee���&V�}�?n� �*�/�N$�T���i+�\,�J�H�.2f�XO~�L�"	^�p�J���B�L�+�����w�O/����̎R]cF�N���}�2HT���8��x�g���:}�0���"�jͿ��˶���M���%�n{]�<$B��<�KK>�f)�Y�*��]Ӹ8��L�F��|,^�'��i0Y��a����ُ
z*i��-�a-���n���6�|���fa����C@f������Z�I�#���<����ebK�+�E��ؿ ��%�4e��[~����p)c��d>�s���l�mZ@ �)K�(:1 �%�%*���M0�4:����~�;b׍G�@��Q�us%��7�ಪ��y;?�8���>žk��>K4�~,��>���Y�ε��y ����"\�A�K�Y��r簾T"�D�d�+����?)
�T�����Y5�}��MY`^D&p�UW�_%�J8�ַ6��Xھ�#"� �:1�L>�#~QRs{�h��T�wXQֵ�@���ܰ��E�<�������r��Xdۦ�/��Q�o+3푆j��7�U�ZcΕ1y�@��i5��B���h�̂c�Qr������ձHE�X?�=S��F���;n�N�@2��Y ����o�\���8�qTzeׂ���uu?e�O�F;��Pz\-l�JQ��7� �O&1n��I���/~�z�bu��玛^�	B�W�(Hрa7&Z������k��?�c����؜x��C=c����|�	�l���ˬ�kCE��3�`ڼ,��/�}��iU��p�.���-�����z
���n�^������n�.��n�����.��CBi��w�����}����9s���;s߲y��X>��ȿط��ю���s�e����\�,T��P(e�T�ރ�Ŧ6��#���1H������Ħ���e���u����	�S��Qj��*�	�7��m�Ɠ�H�ե��^u\\IBhh�$(-�Aȵ�f�Q0$0Lu�J[Gb���e�(���Y�OX(wMy���C�FQ���<\j�ޫ�
������#��g9uM�2P\�7�$���l���&8��a%Ұ9G\i!���1��4=8<M��D�sG�R.$8�t�i��?O		���{�)5�A��!i!�+|cw
W(+:d~h���'̵���X����8)�]�H,��f9C�%�c�z���CF��"V���ĊەC~�E"�Q���j�Mi�B
����ZS1j
vn����&��YHL��y�H�R�#�5�������a��8�߉���l�~�+�YT�w�?�`��;�-�[ڨ�=��[H����M��	e<p�J���I\�V�T�IN��+�G�NPʏ3�_�6��ް��&�C��4����l�;�)$�@\=z�,x70�{�d�|��즨�<lyg�D�ж�����gBi%����&4t/��-�NH��i�~?���y����.�b&��Y]T W5���B{�zGL	���`T���{����F�Wخ�9{��Ӻ���t���|���{v�e��$M�4 }d$J3v#Bxn�C�i �pG�����p)���{��3a�_���.�|]T��5
*�I�{���@��!fo��p���>���l�C�_�Ptq�P�D�Y�`�a�Du��s�����8T� ��:�	h�����\> ��/P��l�xh��s�W.L��ў�j���ޕ_m��6���+Wb=�ڰ�l_,*u3��W��C��Ζ�q�:�M��W�c��\�>�	��q��H+N��7C&
�NR�Y�������()������
ҍ�� � X)����&#^����Azr_2��_M��!_�a>ሃ��k>������Q�Im	�imD�v.��:H/�Ɠ~�m�7�Ó�$�%��Y�o���(l����p�Ψ�1m1�����n�oG��$$�aK����&�ew�o3x���ʊ��FGX�:��2�(l�j���p�1C���4�&�P+�eZ6:{�vpw8�pD�
#���P�SQJx�����G���q���͓^�3��Eo,���s�Ϩ� K�&9J�04���yJ�h-�v@���P�����TCoͨr8��%�T��c�_W�Uz`���o����O6HW�+��Н/}!��7��5h���{ 7�'E?�v�F/���K���A�ra���(a�$fx`�ġӨ�C����Of~�䄧�DG�
�R��?i����p-u���G�C�"��/6�u�X�A��\�	����  ^����-��	T�v��
_p4�<yk3a�7ü2͜��:��섕�Ge�"�l���8"w2N��|�yb��e������g���2~�6αv?k1�~<�������ƀw#6�[�E� ��F��F �Eڂ=B�@���_p��\��^�ƫ�zDǺ!�fK"�\�^��/7e�vA��WzD�,:\�����C_#jk��F#	T�QX����汃H�̉�i��2�-��n�����%��<�����O�9+a�w'�߿G�Fي�%MH�_�:��*��UT�ڄn���Ʀ�e�x�LD0�?�E�����&��5����#zf1bqf�ۥC3�-v$/۷�ùW�~wbz�^��Y�~���|#���FX����oɺ��PYH��O��6��|���6�	�DnVW��!>"^��m�9/Xg��τ&d��*��FKD��G�Y�g��#E"� ����� �#Vٓ �=�{�h �����B~��GL�1�
����*& {��@ 4��B�����:%1�`���x!�	��k�~��:���,� �M��(B�������q
0�����c���]��L�ڈ�L3! � �7��׌��ЁvY��x���7G�$��dX�@����Ƙ���]	���2�C1�\ ى��i`僀|	��(`���`,����� ��kC`?���<��_�=��8 >��?rQ �HC�9�L�_3�L4���杋�� ���@�=���SDv1v2���Ձ��F��y���|��}�O���c�ՁG�z����{>LsMD8<D7�L7(ژ�<p%�,7���p�D����fi�@֩�7��\rB�;8�J���R��U6ǇX�6M��T��&����da\�PO�#A|A�A�m�Z};�$��	���Y�;�}J�O&gI�r%���yB$۷."�X�(�c]0�(v�"�3be�1��u\����P��T��$�Y����xu���(�ڍ,sM���X�b*>O�qGv 8x[PR]��f\�`)Pg��6���el�a�򠗭��Z�(*����g{*v�ct���$y�"Ui1j����H�"���zH�'���td��oHL�#䃴9��^&@9��~쿏�NC��RG=��Y8����$�@@��m�T���%0� ���$G�^0w+aC�#$������ט`�g$�L���Ag�t۱��06��^�����֩\�0�G���R��)ZfΘC�<(��}Z20���8��i	�9�ؖY �m�����7�~Z��x��ե
s42w��B&	��J�Y8�ޙ��:��F/nǬ�2~��ᩰ5�d50�Ӥ�2���S��W�d�zش_ْW�@�����9��Yz���G�T�ғuhm�a��+�6���wB��9����20
�A�� M]����Fa�X
@�~0I�{<�۴���)��|��-X��n,���߯�0	T�4i:���)Af�{��#�LZW���;�����z�;�K�Z��y�p��R��A�1O��GK���ɹ[ۨ��%eZX.�n%+D
O<�\��F ���?�'AKIɏ]Ϟ�w	�ƢN<Uj$�����F�C���������U2e�T"���5��+Čp��y@�k\<l!�mt����_[Y�c�Ld���B��RvN����Ǒ��m{��lbIJ��&�8�\j�2���	�|��R^0��B�'�JBNG���(�.���ç_��L <� ��b�R!qh_��yD��4)!�s�(����W�G������eպ��/<\
����,.$��W���
��ݍ�rI�u���c�Tn���4�����*7�]"�W�%ͳz�������gZE��� �P�&->B%��Q����Į����9�x��=�r�:��7��M��w*	�ˑ�g5R�uEy��tk��)���%�ؾ�˘�yғX�\+��Y��? ���N0
�)f~QH���.�	bs�_��Z��2�5ս7���V��výNr�Z��h}@S���ߋNe�q�6X?NmT����m��m����ѹ��_#�v�$�U� ��~��j_��H�\0��@��"<li��ț�l�n���AZ�QRJJy$�9F��Ht,�����H���o5��kfb���2W�'x��;�1=?�0�KN��+�����c��;sXWQ	G�"��4c�����
A�,۲خ߳W�9�Uq�W;s*�XA�,v�_M��i�2�_�/�[7��v�HKKW�yy�|Kx�+Ǿdm>�k�_��z�1�D�*Ll5�>C�Q=�"�D�emP.�X��]����qǥN�<��ieE��J^ş����vn��iU��}�g|�'�ڴ��	��\��KP= ���~�Hy���1om=��$V�㝟x�t��^b�a��&(Q;3�5X��6�d_���ǣ��S������a����@��գ�n���ބ�adm�#�|��PmP�n�f��T����TXu�y�u�U����_�&ݾ~r��\Y[/�~����Uj��ū<X&|k@6���3 v�ga�[O�xz���F��3����?�2���/��u�O%W�?������0ޫ�*A�u0>�H�1ޛ�%���OnS�qMfHH�(�$�k��w2��+��7��CDȤW'5�\���ޛ����ʩUg�įo`a�F1{�r���R�
���!O2���]�v�� ;�h���꣞��ХAX����5C��q�l(��8���j��6%@� �E�US5��M�R���	�]�]0���G9q�����)�=��G��C'��N��"�[�I�A?O%֭���2Н�����糍�_YPy����v|~7�Bf����,֯_�q�|��>�Lxh��l��Pm�,��Hx'}��W\|��r�=u������:*��<5}��Z=�;O���/�:��KU��g[���7\k$�o3e��X�_�(�\MS4�q����usg��M�nGG���%x7-_�]�O�U�Zĉ���v�X�Y4��-����@�Iŧ���w��o�Ec~�'�6V�E�wE+t[�P�##qJhj��^Sm��>�i�_�e���U���J�v���F;��%�����M겧�|���3��Mh��r65���v�g��4�4���vn��kIs���'噿�t�1�=�����2�xj�ٶѲ�M}@�L�+��	6�5�-c�f.m��f{��}F���'�򢜹r����z�F�~[��������g,U6'��S�H��l��Vos����%G$�6eH|�{{ζ(9qT�H�R]�i��b��YAަ����lXϤ�2I�NѶ���QӷQ�*:���n������0F2?��>�>�!��ԿY�Q����j��3I����֑����	_��댏���5�Ŧ�ٰ��f�@��j3�|͕���rX�0�3��������Z��*o�J��i������Pi��C9j�(8z��hT4-�J'%��O�,l�;��]�`�f�()�;�f��l]��������@j5�U8�w֢���}ޡ�<~H�	�T8]]�4|�1x[�ت�fp��
����m%(͌�R�vxr����_P�!+M�5k1��s���Ό�4���EcK�Ϙ����ٸ��R��>�m���6:б$�Z�� �Rz��7�v͍��8��p�]f�}wδ,F��@��T(^}�;�/q�j�O䝮�+���`�&��D�0*m՝�E�+4f=zH�\�,1e΢qG���st~^	C1�;�q���'������e#[��ơ�w�J֩�����m�p�Y�~Z�¢��O�5*�Ҷi���b�39n��\��]2!�I"��g��q�����?Ȉ Y���&�/q[1���ϣfM7��>=%�w����]����x�5d�`�3�AtC���﫷kMM�hGɑ,z�2W�辣>��!�^��*�[���&
A2�z}[HM�]�I��������h��ao��|��՛��aC�F8�����dɈ�
u=ej]&!/��I�~j~ɬ�m,�f�B�̇�8ң��Y�6<��7/�ۭZ��v`Nc�����yQ��Q`@�ڵ~G
���e,a����O���2����D�*��4���,Xw�z#_�s���ڝ��v��;=�ӶF6��-��ua+C_�� j�'6[�z���S����~�M�'���cg�Cxwoh��P���x�&S��U�\��7��Ļ�����6{��q,%�Z)���j�C1�y��&��T��&	�M��F^�r;m%��jg�O�@��D�8^7]�~�¯�������_}f]�����)XF�p�U-V+.�d�U���6�{L�WC����8��N���w;t�v�m>��s��WV�|�>�y�m�N��Hr�1��߫9`�S���U�d#��C6d25�a���`禡Jq�[��T�f�;��]WǨi���+�a��ɡ�'YY8)c����r�R�ۉyh����=���_o3bͻ�KI�#��ݿ�g����?�Y��t.n����N���0n��[\G����UC�ۄ� ���z�".&,N�"�2&%K�ޖ���G��p\O�g��흴׾�E�@�<R�վ���Iemd[�������mY1,y&<Q�{%l|�t��V����G��F����5�l7����H�7�J�GsӶC���lDkd�q��y_@���T���?b������g1D�~��6Xq�vV5�aI΃���c�������C�d��n�n➦��n�Wn�K��;���^���ܤ�9�㜏}qK.��y������x��b��j
���J�Y	����[�ͭ�2�>�BR�)��Kҋv���B$����I�k��� %����?�qЕ���^'YӘӾ�@e�KN?�#]���ڨ��R��'����ϵL��f���J�7����ܙ�Ÿ� wL�P�7� �{��C$
yLGP��1 }��

ڈF� �/
5�Y����R�j��
���EI��;��x�'̵�xO�W_5��@�K��ymn������z&ju���-�/�Y�<|TK�3.7J���Ê�Y�$���UJ������]���ى�Q�I�+�1��o�I�p�rz�Dj�n߁�����RPk��ت'x�+�\���fo�gG������[vxʴ�O�Jc��!΃��Eu����K�ndUrR�
��Y����C�h�#����樓c��ܻ�@R��%pzn/Fܶ����=�=7��� ���!�����dU��s#�=�aA�~�הå���
��_�9'�TM��vfڲH�#���\ҶŲ��gB ������
�XP�[I>����]�E~�v����;�315)�YY�R�C���x��?���a�Μ�Z����go`��TЦ"E;c}k����p��A��5�1�Q!�Di�B�u�op�8}��=^����uO*�����{.���8��$+��{?[�]��s톇o%L�ޔW��P��"a�����)-�B���]l��V|Lq�{⟤�g��V~+>=���o6:4��t
��T(������[��R{R�8��ɻ�5OZ�8f�r��7��d�W��xb�H,4���84]��ܷ�䐃!�=;�����	^o�FL�#�5xE��x!����m������]�����IGo���s���%���n�*z�F������qo��NDG� 1BG<z�skA)N���i/%�oy����:ُf�Q�׿���2Jw��m[���J>��uD9l�F��X�ٸD���I�)j�D����C��#!�_������zؖ��HB�*Z>{��9È=��A��8/j�jc�؝���H����c��,��P���A��g��j�v��
)�l,�����+&(h~��~w�����:X\�J|�$���N�l���d*�����9iV�$q�i�⓪9)�&ڵ��9�	�ߖ+�,�4�J�4,�^��u��sf~!��o{54�ƣ�dMv>�R�$�����a�@~3�A#g�Ol-�l�~�R�Xe�3I�x���s����@�M�\8�(�:���&hH������X��<��PR*`���ӧ({ *|;S�H�H#�X�7�	_ ���mS)�-�m��āg���b�"k���g��3㧣S0�m��j8���F��~Z�h�Ż���fC��3�ë�E�$���������fo.+�'s#�ȉΥ�Ѳ#�%n9���X����2#�S�O����s=�|�j���7q&$�F��6�����w�8(�;�e���e�Z���@�r)�oo�Mrko7�g�Na����_��!�G~7��{��F(�\��or�|��z�p�Ug�T��Pdq�ט˲��e�����u~��Q��ޫ{w�G|��@w�
8L��x�����B���Ƿ�͹Zt��mu�+�_6����eĄT�4��Y(�YNpHX0�\��d��N��\��"��qk�b�n������ڈ�x����/Ls�z4"x��_�Y��D�n����aj��.����Gb��(����L�["�v��c���G��K6��!H�*FIs�������������W��Dl��1 DT�����L��z�T��=_K<,Fg�e ��
�d�td3���y���W&��|��0����o���9�YǙ�fC�ȇ��-�Û"P��NG+�O�\�u�O-@*�r�v�"�⃃;de>r�k��q�i1��jI[W���(b��xE�Zf��l�g�??;zFR��'n��pt�y�z�O��=k�AGl�U)���]'X���8Q_0}g��%����n?��:c��$Fw{X���{��یVDn���)fw�>�]��;��3��Z؝W�.��I�OɋB��M	�u��:ݖ����:.��!�MBP�]P;DI��y�ʫA؛�!I�G(*��4�ȷ�2nn6�P��P����堁Gp"&f�E� �������oE��g��9U����0�����������%� �i�ȕ� dR�p0<U�/Oi���P41�����5�7[���SL©7k؀ur��Vq��h�����e���,'C$�
�qC�?>m�T�)�`
��P���fٽMsa�Y��Fq/p��Q�չ�\P�I7�@�!�#�,�Z������|�BZ�r�M}�FΞ��{Td'��!�ԙҝk!�j3��>8Q�	Bw�nq����#��v��yjpؑq �h$]/ �L	�RЛ�M���]a�c�766��-Q��#$�]Ӳ�כ���:��O�D�*=���(lU-Z��f��P�:#����6���
����w�Y�W�f������Ê��8 ��5�ݜ[���~y�&q��  ��m�P��q�R~&��/�p ��/Z�����]�4�Q�TD. ?��~jU_ۚe�gi��ݮ�Z$j�hh`~��rkG�4d�	�)n
���-��모 �w�t�r&�gqo��<�p0d��q�S��i!��g@��	/~ՓRٺ�����f���fz��$л�m�
���|�9Aշ���OO�7�O;/&�NO'��[�c��j�����ȧJ͆�Y݌iU���:WR%^����`t?����vW���@�9{׀ϥ7����~�r؛w9L$h�C���.G�Զ��翃8�t��WT��;���ά昖�Q�a�4Й?K��lji���&�vS8`��$]�^�������/�k��}Mޯ�+�}}x`6�y��]��śY�L���
y�b�4H"=wL#yq��-�����zI�����w��)j(`^%^YM�;��k?H�#`�h^ȴ��z�Q�mL6�!�ޮ�x�6���~5���n�o�>���d-WQ��@?��[��2ş�o.��c�vB�J�k���Q����g�����3Y ��&��!���+�¦⽑1!C�2�؈ٿH!�ԄQ�Q�)���&t$�q;\�Hrl�B��\��J}X�B%2�>�H.^�������M�ڃ��Pb�2��V�ـ��fYԆ�u�]�냮C"B���N�8Q�!iTu)
r�1�Ȃ���%���`�"��V��}YP�H.�ʗ��7R?�=Φ�����^~)@���)�i��	H��moy�;aW�Ν�l@�t��`H�����5�����"2$�']JE�!�c]�.���zs,ܷ-��(X�nr��+ Y��A�M MQ0�6xYM���r�5���7�3�Pfn�=��T��y1��.�7��d�:@�{h|������8O���g#ٟ]�╡&;�x�v�-���[��)��B��gRj_ޜ�i�^!/-`	���h�вe�j��J&A���3XE��%Ƈal@��H8�6��t�YJ����Y��b�f(���,{�ό�t�)���x���:�����y-�%cz��n/2J
��2���l���4�g���$�,���a�J�G���Mޔui\f�����������?�a�����97&gi:Z=՜#��
_��]�;m��ځ�[����_�V�$.k� r?����srw8���ڲb^㊚tɋ�� ��qj�^l�yڒ���>��P:J���Yo�l�?��}1^�f�s�����;��w�� �W��*��W����ï`���m�C�����j�-_�?԰a9��@������N��i#ˁӄ�.��l[�g�^��:�n/���$έ�(hJ6n��؈��v�5a}��&"�g��9Q������)N��y#��:�y���Ȫ�����z��{����fUT���l�����:���獉x�{L�ʴ�d̔��On�c���Z7���s��N��r�	��Yǆ7�pȟP�o��-S�Y��>
���Y����& w�5�Z�~qI6|�6ے��ъR'f�1�ϊB�~R}�v!3�����N�?_o|xIm
p�0!��$���	�g�\0@S(L���1	�s�{�`B��-��^�s5��GK��f�Am���+>�?{\�d:����ل}�78�E�X<B�H�U����0yE@JJZ�٬�#�̌�M���(����P������yO��y��oK�l��2�˦5�"��b�L� ���ojh�uk߭fu�Ƣ�4������J�U�k�珙�Z��M�\Q�z-6D���za�:��W�>���N�8�_a�[�����uhE�d����m �q6-��P����'�F>1m/���?���;�b�i�fy�ۀ������^�(f�� ��{��n2������0%ox]�̙�]�ޏg��`�yv�O��~�̟k��@�|�z�.9����2���U�w버�vۚF����q������+j7+Q�-`=<�:q����7�SXpd>>�H>n�Ds�
��*�}inv=�GVB~x�I�K5L��,(e�%Ԓ`X7W�*�x���ԗ�`G^���u�J�Ro�Y�H*�.�")��k�۽Wm��Z���/�vI���-o��4���ޛ��_W2Rn�E��� ��sv�����/^E-��rȅ\��4V�s���u$�q���>~���8z�[hr2V�E�]�U��N�l��癭$��c-v�R�/���Uhl��y)bxnW�n��e.���`��L@���{'���+�T��zye���:�LT�J\��]^6�&D5��
q��?*�w�R4�WmY�o��oߟ���A� �n����M^�-���7nhw!u��
�4��7"���V{x�u�����#B����1c��G�e���+�\���!�8�.�˨�����d��֦,�j��j��>d|��1�$�T������b6����k�(u0,(�/	�MB��N����T3���h�u�CB�g�˞9�B�'K��l9N�$�M����b������Z�ga���*��b�HH��4��@gͧ�ݏ��n^Ϋ$�%~��U�Ȁ�����X�4�i6?B(��Zu�8��Rw��'#��߆�L��Y�i�閍;QR�6s|�)́9$� ��B��q<_��#��|a\�#����Q	\$N��=j^����H��z�Mrˀ�y�Z�V�C��QeU�2�Sz���#"���s��i�2;�e�w��e�^��">�8h�62�̅�%X�?޼�V��Q�=]i��]o�=�S�gI�/c�oX�q"Ǻ�mr.�/�rq���>�s�ػ[9�_���)[m�rg^bURiE�Km)r�S�Jn�9f:*!2HÆyf�N�S8�X;��j�)]e�S��Hz���g�[^t�#X�tq�9�Y�q�p�s�����U��y��J2�n`j����c5e"�"�n`����>�R�����\��tg-&QՋ�6��V|����������t�b4Z�f���$�����"<8���8E�$���0�l�mڧ�#|b�*>qV/�����f����J�u���.�����D�<�7$�D��<��t6�+���T�9�8�6�'�������"�f�ń|ؿ�,ȷz'�Ũ��3#�����k"��b�%���xN����n��-�lL��&�[fg)Q��K�4tBc�ִ���{B,��5O���͟��X�6��U�-�����<������ރ,m��I4(�GX����󡤊d�-t�8&
W�o�M�y΂B_Ү��.dYZSd���d�׵����rF(3o7�����WS��x���O/˚X��ұ3�����TA��B�u�?��>�]��(0$�y:l>�	*(���v�a�t$�v}B� ��x�!�v�΀��Nm�w�7�={�}���v�n�m�	�#r#�y��`P���}&���Ԭ/����u!,HRlX?�y�h|��\�h�1�w�֍!EAN"uv���]��C�y��$r�~0z:G���<nD���|n$�CՋ�&�r�Nԝ���8��yP4��<A�❎_W苾��7��Ⱦ�����?c���gz|j���ɲ����!D�d-���.�hF��x7�󡯹GJ84uF�ɥM)Lbj�-!�B�ǈ��8V�ܿ��%3���=6�O��x3�⵿D��ў/�1�Agd�EDm�8�f�/�޾����OE5��o�}�adv�ԗ�斾��'�D�v�VɴH�"��"-��s�kܘ~x����X�#�"}d.Y�;Dx󼤕m�-�_�n�GK��x��������߶��&H�{{�4�k�j4�pr�Է�-A��>����{������oÜ���x�G��2c1����p��4�]Ь����`��]T���z��~�fQg�(e�x6�M��I�=hgH(�]�'�?f���=.�[�H�g��/�h�)�,�|1I�6�d	L��!�zt�������@��Mh��ʟc��ҵ�m[�s�SH����|��f� q�d�pU�~�w�r����w3�e��YI��R�r�=ٱDH���kC��Fl��y�w���3]���B`M�����h���#�E��H������n8��`퐲
�K�n�EU��5ii\0�$��%�Md��Ekl���!<�E��1��[޻�iB�)�e�t�}�������{S�@��0��0�d�yQj�S���䟃01��m�K��U)\sB��ŦMxBG0�1
H���&J	>�q�f[P�f1���@1QrX��2����գ��Q��O�D���s\���L!j5'�Y�D`����g� �0�8l;��
"��96�)�A�x2d:)Da��R�,c�{Q���JJJ�@�',E�$��̚$P�c��t�^��T�2�%%���c �B�sCxE7�?1������YD#PL���|���>���͠% ��'�GH!z$A��_�L \F��@q	�Å��B��,���i$�OC�� ��A l��DY��� ��1dL=v�)UȘ�a�7�Gm�cF�멂B�2&��y���<d��;��� hMA�cԐ��@O~@$���(�_ � # �2?��	� \ ��Lq�z�\l���	��-�ƀ���`˷@hH���ɮ�TK A����_�V����d���qBHH�����^�
Ї�	�U�7��� �4B�O|e���} nVA�G]".7B�&� n8E�`��-NY��9�"ȍR�jV�Y�X04�/
w�B0��C���� W��}k}���G.LKu������J��ݚJZ����\�Aue�\D;j���ҍ�n,}�He��
�su]P�����R�֒�y�z����K4D; f�hp2f�U���n�J(��t���!�ȡ�ЬGXE���a<��|>kŏW���%�Wt 8Z�� =J"�%�ݖe
�֢ʐ������@�]��z�p�}�9W�<�II{���eL�:p�)�Yc�z�)o8�PL+顇���>�ô���j���������3<�0�1X�#=��q� <���ML+�����a����ĢD�oH��F���u=���@�A���ւ�B%����p��С�N_��Q��ç~���MAe)z\H�T�Ѫ�|W��LA�2h�ܲAl0���;1�nO��%������z�0����RZ���C�d�Jf�O�[5�����.y� 0�̓������. u�OH���ej����#��J�<w��&%>X"њ�{��f�.�%A��H�׃5&$�2M�K���	M�
�#��Ats�Ε������=Е:�+�E�"D@�����YDm�����u�"}�~nyv�VZ1� �$�VLF&�2�R�6</�Ĺ��?�CaN'��}G�̈́����CH+�m�+�X�9����`��\I-���n�C?���B��p��s��Fɰ��'��������ԗ{��=��j�Ik��%3J�mw�]I�bO6���C�V��&B�� Z0��6{���|c$�4%l���=#�2	�9�F@]#,KQ4a��A�[�����x�;��Sk���䖂�Z�T5�u����[)"��2v��wA����[����?P`3J(㨈H%99Bz_��\����b�,�v"L?��D(L]$T��^H��0�a(�55�0����J�JN�8Jəz�!���Mͺ�Q�!۫u�4?�k�� F�%,���,	���/8})N�o2Wc�eպ��̷o�۪)�NK�wte������d����3��R@�i�:ޝ���z�TdrX��Z(�Bd��g��	���P޸=�:`�Y_0�!BOa��X��Hsr�z�)�u
,��(0/-)�v�z|�v��]d1�ߥg�i������ć�דɝ�
tb뜾�%�v���<����zT���PW}	�3�,�{hx/�=��$D�׼�<�z$"�Ӫ��.��`.����2�&���K���C���Nw�2�m�J+_n�%
dͽ��J�φ�)y1g�������:�m"�b'�L�pU҄���@���7��w8�� �0`P��(�����m,����>sl��;�ii�Hʭk�FKNr80ڜ3`�;{�E��s���i9��~^آ�GC9p�?�r7���#�
���I��K�i~[��4,�����0��`9}`���c���eE?�a9O#W�Y� =�f��с�-U������M��@��z�G������8���.F�?$ӿs�C�/��ԉ�6�j@�V[;�����	�A/(�O)/�B޻��+0'��u%8lG�`70vk}G
͂gi�%=��B^q<Yn�����'\Ee���םߴ�:�ۜ ������.C�^ڣ��k�tf�B���<s�n�W������ܻ[��n�͏c(�\푩{��]��zm�ٷ�6W��w{�y:���УPJJ. �����RV�g���У����̛�O�]CԳ"�vO��?���`�� �3=%I����@ޭ�D�uE&�����o\?W��=�ʳ���My�z��3����4K���g_ֿ=t��i��7��j��
v���������w��0����F�Ni9V�N�ibF7	��h�=[��~��M��z�tzZwv�����Q���dK�z(�l"`<p3�+�y2��_Z�����e�&j� �"�t�9W�\c�c���"��-�Xi�F��Vp_ֳ�\��rdL�r����;.��7�0S'�DO��E.
���EW���zsa\�����OnE��J�*#
�*8���B���DU�Ye�[Rum�FS�v;�Ы��
s۽�|�^��/�YIH+1]���5���Un'�+_/��U�	������|�K��rr��Vh1��VQ�f�D�Ƶo�6�x[︓�x��#"��5o����ѓ4��I�(�	lc�|&�����x���m�׹���c���S��8ΟK���{C�^iԹ��\a�����WN`��<|���&}��ix��(_}��*%}w�\ܳ��'X�J�h��R^�:�k�뼞�E����wk�ظU���x7��sy#�	]4.�V��t�G&�?0���㥿�7�;�8��R}<�(�&��;BMh(��A�K\Ҍ�x��B�:�5����d3Ld��U����w	^��H���>^v�v'i�}q"�sSl���Q�����t戻`��
+�����㺂��j��Dna�ͪ��D$Y�l�E�o(\&���a�\�?CJ���	+*��頱7�"~<|��:���o�'x�ƭ��ة���>?P�i�V��9��uP��ww5l ���6��"��1�r���Ź�����3�R��V��u}
��<&²(\@K�_L�>��2�I\wҶj�Ĺ�J
��#탡gSBjF�ƒ��
k���#���7�x�����FOQ���g
�?���:ck4��������Fz��o)�1;-;���*�[��?5 ���Mit\d���Ģ⇗�д��_<��+Q�ZQ64��Mւ��e�R��W�*���?^�^��DP�E",�̭.��u;���R�U��
?F�AVn4u?f�����^������>�P�_F���/��q�d�m�4�,��h��{qy�˾y�h�IP�?m~J|"y;p��$�R���F2�h���%��ػ�}����-EG� �E?��l�	���M�C��΄,yL��4�g���}��5�8�?C��.��p��٫4�mQW��,��
=	�һ6�e��H���x,g�:���.fs��@J�(���8\ǷĆT`h��n����t�w��f]��6��@�������$��,����}I,����j���66�P���k]{i�y�oI\��*&��Hd�O�Q�:&�D������7���YC(R���
Fwy���1=v4V�|˪����������i֋�Cpw'wנ	��N� ��[p]48�eC�8���w�9��StwuM�SO�T�HHĊ�IdE@H�Y,��[\�� ��o1�x�U�AxÜ$��i�݂V�%��SC�	"`t��e���9�D�x����!��F�d�������8smK�XWE����5Ua��i��Q��K�4���x��qS�Y�q󩡀�XP��Z�V>`]@}��Dx��D��v� ��l4P(po�o� �x�6ɁE�����{y�<jZ����mxR�-n����������*�rg��(��V�y^(<q���J��h��u[�,��V��ŗ_(=�hv�d���r����7�%0rW\�~��72jʱX�f� ����].*�m�2Э߉���s����:�����3��<W�#dsDX��⌬(Y}�[�6,xb�NM�%�̻첎���jyJ�]�2�iw��|l�hx�\�s�ò��b��45��9�*�p7ћ�yR��U衭��C��<&5_��)�	��x���rb���{s^�u��Y�ga�F�u[*Cr!�r��� h'tK��R*H��go�t��V�E�z�ѓF��=�7�w�R���o�UٌzL^�?��K��(n���;:�\i�4"t-�4x5֑_|��MX<�׿`Մ�}�G{"�r˶��������z��2q�^���?��f���|��G���Sr�s��&_����d�Z��2�_��]� &��w*Z�r%[s���a��(}�Z��gVF˦I��ܲ:���#�Z'>����dv�w�)��]��	�)tb�<+Րe�=�vվI���妎b���H�<v�7����/�z<:Q�?�q��M:]����u���ʴ�T��΅MR �<2v�/�J�@8��]D:�Q��%2gh�:}�,�i��9���o�/!�dwYV���^q�
�Ԋ-�m�&dl��r����뉤�*�U��6�b�M��]�y�1=�$�b����t�w��I��c�ȤR�C_�`_�ٖ�O�=yqa?޵��)�q��9����6X�|,ϸ�'0X2ϴ��H��2{�V���(��3$��s�*��/�q��#U?��@�ɋՃs�'C��/}�6���{��F�G�ۏ�\���i֡�Xb��{H����|���k%}�֝,7��`��-dI�-z'�8�:am���zE�Ǥ1�hڹ4'\7���+U^}�j�r��@*$����n$P�N�-�!p�ϩ®��l����r�Ѡ��r���@?�C�x�C{��v��K"��^G��N�WN݀�������51H�K��K�����e\i�NǺC o;�/�d�u����%/������(�r;��`���//���c�A1J��/n��P#."��h��~�H��"N4\veÆZl̘���!�� m�4,��K�j�G�iR!����۫=�'u�`'��&kt])mM�Fz��9��'W:�OB5?�����ƿ���ǘ��3.����������n*q|ij�fp�w#��*NC$�v��g�>�i�����_��<xT�t ��<K%�6��&�ƥ>FW�9 ѢЋ"�f�|Vwx�ơa�h��j����l`����[u5�<�R{3�-+������!�����)J/}���02.� �4���m��h��ލ���J�|Q�aw3�u�K���ɠ��\��կ� ّxPIG�PF�U�jd�,��rļ|��C?��í�צ�i��H����+p�џ̂�����#+T�
��N�z_���U/���#,��dQ��@��Kd��Ih��8�	��
��#w���2���H���x􍖟u�9BPCC4u����ۡ���B����1����n�{�Ȋ} �J ��L��eE�'RȖh"�/˙@owp�=��[��c]V����휾�V�R*���~��Y��S�]v��k;���e��*z��h�̞7�!&���X�Y^�	u��KP_�Y��0P�7@z��$�oC8���ғz&7RW=� �F|ƾ@�\>zq7q�J�b�dtՌ��](K�m/�����G!Z��U|�.�>��(}��~����
�)wp3H�2l��F����x>T�����5�<DJliYm�So�̭H�" ۦ:�j��t$�a���$V�Q'������|8���5���$����g����m���W3�XBlы;���O�庋�(C��H ���"�;�8������{ON�Y{��v�{�ͨ�
��P9)a �B"aO;%6ؾF�I���ʷ,�.s[��ǚBb2Q_�J �����[&���-�?=JP�/Z����o4��~_�(/����;b�L�U����I�ʝ"R�{"��d� �'ר��� �V���[e*W|P�eQ�ѩDve ��>=�!���m1��bd%R���a�����(�_ZI���?qб1E�d�.���Q��Z캨o�`NQ�NX���)A�l�w"H�Z���b��A�[��k���n�Z-��|4��
���,h��h3���&�j��|�������o��@Y�RqH�2葺�����}��`�c��-տ�Ge�n:�H����e��"�V�%J:J��B�=��i6�*"�7B�ą������6bg�6D��.��*rn��!��Х;bI!Գ�����B�X��jK3ʊ@���O,�)��/}(�7

��,�6�Za��Ҷ��7�E٭����k��Gm@\tZT�_���%F���┯��^%w�'��B���2�g�!�3���[Y5���a(1`��Ƕ��~`�uG�@���Q7!Ͻ���g"+z������F����I�?����T�P^B�G�A�W�����9����~��DcΩqB�O��z�w&:ss�d� ®z�t��3����Rm�ҽ��w�����nr��hy�"2B��Ӷ���ِtRR�mv�+�tY'�_=7L;�	vh��N��!��+�:X��'A���;���..�W(�j�5�Z1c��t��v�%�p�Ә�M��#��\@�|���/rW'��f�F,�[{�Ȳ�~���r����6Q�x윗�(�KPV�;TbJ�<$��jW�]X ֈ7�X��������,�R?N%C����E�`R
�܌���ju��	� �i�;Mo
V[�j�C��DS�@�+D �9�꿛�eN��n���q��_sI1�4+8����\��t
�x~��hyd���3�L�wE�l� S�1#q��"��������P�bd=���Q��;N1(�-�2_����b:
47��v[�;\��b�^��&�*;6]��{k^z�qл���]������{P��ǥ4)J�w܇�TS8&�ʴ����e*_O����4�N���΀%+�7z�)J��Y�ĨP �Q�X�����Y�7�c�\5d/�&9z_��b���	�of��p�O���O�9)�Id���1����(��{�ח#E��Of)F_.?���t�҅�c�"�t��{B�H�q�[�4+"#E��;���h�l-Ռ뚮��o�sM%ay�Q	�O_�~�oƄZ�
]!����!��[��z�*o�m�z����0��hL��V���_�yU9 D���ߧ�_�Ї׍���ޜL��Gα�[�>�˲o��HyC}�k}5��zuB!����rQ_�AR�wOY�26}�;�B�c)��������K,��0�3�̇���>�=��h��t�s�A����,	�u�<e"�l8��*����rP@�ظL*�y�X�,P}��mCF��^R�Y���x�j]��x>ˇ��wn%��l�ޛ�bq�4�[�����Z����~~*ri����{�7|�!�~�)�m~(���6��]�eHS�S� 4�-6�����V�E����.����5�+r��R~���1�9��lF�(Q�1��?��J� �IF�tJ�O�Jz�oO�ǡ�c7���r��P��B*��60�v��86��*`�J(�����T��y�S��@��y�m%As�i#��>��\�84z���:��ڷ̯�[����R����U�Uk+���ͫ��,`�g�"!/rF��.�u#���DYY^�?��ӱ�K�?k�� 4�D�=J�_���+�|Cy��{D9D�?��-���tQΗ���É�1������LQ�%z�K���OTWW_��tM�8�"��T��^{ۘ���ϥ�p�j���[D��y��@�_!HD=�B�ᯁ�)t��_C�V<��V{��dr�H�q���vλ<	~����epK�t0��INN/�Ȓ�{�7{d(b�}�]e��;��(�33��j�(�~2�����V�f�+rk�ާ7�'+2�����b�Ic��R..G��y�ngG"XKR75�p�ku�����&(��qSJW����ɚ�1M���Z�	���'X����{o��ߔm2�$��B��F������o_�A����x/���˟3�䥧Ӊ�>��r���@gBkΐ&���,�d~,&+xP<�5�ʹx�n������p�i܀�X�n���Yz�K')�(U0�����\�J����_�J=�Ʉ,їǕ�#�J"�N]j���L�����|����?Zdu�H*�U��{[8y`V�~
����a�y�Ƕ��(H;9�7�堣����YH�� .� ������S����ղi�W|O�8F���_l!���U�L ���b��i���b[_���Ͷtʻ�R������B%(�mn��I����c��ؚ�[,EZ����cf�>��SRRr�U�.�3q�'E>ί��=���U0��J}"��x�U\�?T�A�M��j׌����o7ye��q|�n�ئR�6��[[�|k�>���}��_�5�K�N�u�v���\V�'W)��5�x+�����^�L����:v~~�$�c�+����B�]�l�mN��}+u�wm"�n��b���qy�Gy!��o���Џ���Շ3p��8�@ɯ*P��q�@2,����f�-�݌u�� ���O���X�`]V��n��O�\��A��c�ҴV�1p��_�/G������xq��`҉��"'1J��r�~��D��C����B���)Uq!�


��?�X2����$z���^�o��"@���Z�/�>lhH"�Y��Y���x6"�y����v�W������'fi���g��m�<��S�8��7�̕�dv;/��c�����}�E6�'�@)�Uw=�;c�*�&��2����� 
��A;�nLʆ��`
�ϛh�������$TT�g�+'�*7�P�H�3����E�<0�#�'B"����=��sN4��fah�Og� ��/����c����:�;��綵�m(��梸wz����Mπ�Q��������������+rr"@��5����ɏ�b���e>����Nc����!	g�2m�:������"�J?�g�%�`�x!�A�÷821s-W��y���>Ƴ'��&�=]�:��f������'hb�l2x�FSs~x��$��V����&W:�֙$��~�E����#q��bv����x����Q>c��m69k�;?z�ld��,ž{~�L���C��)J/�v��a9]�Y��§*m�!u�z0TI$/����!����廁���"8�ը���;�$r�/�!�L��i�8҄�v�Z�!�XKk	�(���"y
l�4�����t��)J����X��P�"xo�iD��͸���h����djf����C9�.����3�}��c��j67�OJ �Z9�!	�H��,X��R������]0A�͙sjt}
K�b���L::\I�4$�*�ڒrwԛA�X�OX��z��Uâ���L9��Li^��Gg	��f�M������XŹ����CJ��ě	6Ĵ�	|:��;���� �c�oht1r����Gw�;��z�+�\�l��H$ܦ�ʬ$H6����<��Y�F�i�+{x������q�5��-�:��>M�J��	�'���Qw�"d�J_��&�����p*�6����u����W�{���)ծ�x9�-Q��U��m��o�k��#�\7]J2��hD�eD�����?��ֽ���C��X�������.���:�;l��}�dU2Ǉ[��oRA��;����\")��`��%4�B�;-�mΙw+Y��B��ze��\�p������H�c+�M���l�u"��Ȼ����w-���N�K��d�_�}k�Ά,!c��`�Q�V�KM�	g�]�.���~�^h��7V����n��z�馁f:�8���v���Z�Owr��{d{�J����Mƕ�G5�����6�s#�U����D�������8�k��8&�p�KWzcޔ�f/��\*[*.ʺԅF6U���ɛ�]�7���u�VD4
O��3���0v�]dh�g�|B׍D�c&�pv�M��đ�u��8@\A��Mb��S$Q��th��AJk���b�E�{�5�2�]����0DZ7�|������z���ߏ(�¶r�D�7��!0���F.���bs�8A��#ѯ��_��
�x��p&V��0�ND"QD���N#�ۏZ"�ʋL(ڷՏ9!V������$�@�q�<bһ�.�_�;R�l�$n���Է��qbuqq�`|z>��a/"��$�p{��#�1H���?��mp}��������v84 ��u5˚�OSiG]����_��eR��;��Y�X0oM��*�6>�U;�뷁��e��b��J���-�k�Zڶ Y,^y���ɫ�A��yL� ���_�߮��vbu;t��,�ݬN}Y������K���ak]�F����fj�A��Q��Nv?�ޓ���_(캗_��+��dmt��b����)>�~�$.r輫*��z]݉������)aˉ�X�)Z�ɣ�s�dc��E��5è�\��?QVģ<��-%�RsM��*^ybȸ9e��U�ü6W�c�D�w������<c���ڄ�$T��������s��C��!�� O�7�y�(m������ZX9k�>���v~�P<:�Vz�B��Z6�r�ȍ��~1". U�M�d19�l���\l7�KRn;�:�f����O'��9%:�&=�;[Y��vd��{n��~$®���x;	s���7q`��؉V��0Q�m�gu�^���?1�5h�ʢa�_��։�Ly�9;ǰ���!����i���^}h�pq2,m"�ɮ7���+������Epں�e�"܀��j{�PC���J>�oz�0X��]8������R�|J��n+r4��F��b>�qgk���k����Ã���@�|�Lx�PB
�wv�iQ�F&D�!p����L��t��U��i�U~h,'@���4��)�x�A�G��E������UV�{9җ��H�~����u�$@ko14�!jY_a�p��ZI*l!־�D��ؠ/f��� �Wg�V"���`�/��j�kz��`�a���
�G�s0p���'â�řR��o"�{��I��)�؇ u�_�Vt=c���?��2߂1��F�D�;&$C���䴻B���(�9�n&)�xs�#9�����?{Oh="_`9f��{"�=E򕇝)g	&������q�|[���{B�wo�/��2�Tžz���< �VF�$�5�.��a|�%e�q�,��Б�i�iB��Z6���5(YKV�����U�׹(À��,�xP+���Z	�q��g���d���T��T2��� �P��X�Tl�Qh�S��%l#�vZ
�u��h*�Jb��X��i~�T��)��G�����{��ϗ�Ϻ#�3�y��*V�ޮo>��T?�p�;��B�q�U�)Y*����9A�����	Ů(dL|��Sr�[���A�G�⛀��&�/���7:��	�*�34��G��*��L�d2���dɘ��p|���ld����Z��{��i�e,���C�2��@<"2T���/XA-_IB"]��k:	��,��)L�&��
�`�$FF2r60\ƄΓ��Kg�O"c_5D�� T��,�ʩu��*Б���E���h,蚜��yp�Xa
1�І�(^:l�f�J�0�L� b��"0�%L9o9 ]1��	��}�9���
tM]蚭�yBp�Ԡ���������[�	���*�Ua�:ѯ���F��D���7�-t�tm��C}`Cx�5�`��-j�E%��HǀjD�Hf�\آY�2��U�#��g�NK�CǦ�G��( f"Oؚ��#qÄv0!t���1��U
�֚*4D��/�*ĀY^U��Y�(��ǍT��b�B k5.\�'845��kvLv��W>����}���Մ�°Vl\NN���x�̆�!Z{�86�Pl,)�e9><��"�"h���p��#D�>��/���uR���Lv��?�Ċm�ɚ�,��JDφ�;���~+��=:>��_���N�*���?T*Ygr}?i��{�E��vme�:T�L��Ǝ/��a��U	��?������P��k��h�P�8T����Ăr>��b��p�T4N�"Ƥ�q~��7Xj%��Hx��%�퐙@�՚k������'vBK�R��6{\��I��q�H�lh�=xı��E4M�+䉛4�,yÝ�
n�#{��"�1��ό�9R)�\��X �j>��i�F0.��9�$J�S:�m��.��n�)�@�}�N�\�ԗV��J1��	)�N ����:K ���s�	]~��/�Jk7�t*�<�
!RBQܲ ��uvb �����;����OLF")�S�M��$��U�,=(�i�_�`�%W�+� �سy���Xٚ~{~�,�vI�<�=@�.⊆	��)���ЯLC�~qi��ǡ�C ����p�K��i���W�)��;���<��8['����C��%t��N-��zMm#��϶Q��MH��2��T<�α�И��Hs�}�	;8q9w�~����ާ<v�����QW�@(�N�w�<M�	Z@����!��l�_�@ri2x(��H�L��ڨ�$$[/��cg��	=��'| �͗����]���8�}�d���y���&>�!F�)�NN'Ԟ ��î��G�R�~�z֘"N:6���6>X�����v�:}
K��������*�D��Bʙƞ�^_��Cz�>�q~���䙄�^��>�ʵ�_Ez� ���z� �P?,2�{O�_혭������70���	7���ށͲ	ox(��;~�� �ꨥ�FQ$Ik��9�~�Җ����% ���;(�a=�Ҽ��0�ɍ�M�����u�[x��<f��])(~�rM*Ǹ�W�2M@��S�G���}P�L�o�+,w%�mu�^
�:c�4��ဏ�?tx�P�J0�v�_v�GD��;���7�x̎]�=�=�>H���[ͺJ�m��
Q��e`!�|�쌍W��H���F��B8�n�Ф�74+m�Y,�'}Z�70
$�6��O�C[�ͤ��r<���A����]�o�9��m��՘'����4�5$j�<�JE��c[J5�M9�oId~b Q���QE�֜]̈́�~-��o��\T]�6�1͕Z[q�b�$�"�=�rw�%"o��P�d]=�עr�~jv]7�i��3Ncr�ӡ&`?2��;�d����h��*W M��a�,Ǩ��om-� �m]��N�!� ;��=��£ܮP�h���� x�p��b�߁��j+��C��+�	�{nP�}(?�Wc��(�e�ɈEL��~��C����1����v��Sf��;u,x��Q?�/�]Q��r�GFPEQ��4R�	5"��	��-�?5TlP������#�G`A�|� 1��P?�w��&o�����@��4�&�5��w����d���K���7�]r��C��?n��w@y=mN'�`o�F��I2ॺv��d�ȁ�O-��\�!,`�GΆ
��v2�㈡�@KE��F���J(B[�\>cTi�R7PR�M��b�U1��bj
]..+�o���Ϸe�W�����z�?YA�Q��i۱��E.�\���1�����G5�+��f$��p�������m�b�����:'���~%%0�Gc��m'|���?W�BL��ʥ����9�v��;�l]���q޷������~�ތ?NO���V�Cى�|�{Z#�e�*{!g&`-u��SI�}M�[�����p	(��d:�wVds�C��%�s��QT;�>H�o������ �^�A���&%��{u5:�LD�)W��Q�K��i�1;���yV-w��&����|�j��J�%��fcM�A(�W/��A&!74��L���޿J�m��^�2�ͳhǢ�O~���{[�(��f�0�.k���ez������e�+�Q��
���Ϫ8���+Ø�G�MNn�Cdyo "�-o�b�ܰuI���u��"L	>s�pI��R6�6��!T-�r'��G�(��ZQ�%3	�vi�li�~|���/v����~I.�*<�r6X�+�s���,Y�v�cȘj%�7g�*"��CG�#��(����@����-�jq�X�ޛң���-���ȷ�.%6���n'P����я~�$�,yM�}�X@� z�s��k?�-C&{ �^QÚb����`wn�|�QN��o߉�u�$�T5�IY"�Q���Mc�}o�W[�`�?��ސm%����h�-�]��hdEt��~K�$��vx��+֎�w+�ް��4��tJ�+��Str���t�F�y�q���C#6rT�@�J�ş$��mΣ�6��>�L�S�D��Q@��9�U�$@�-�v�cJC,*u���fۧg3
�(��;�.Ń>��z���$�x�gW���[9Ky��1f��o�{���b~����;��%	��X=���Ka<N��D�.h��#���y�ļ����^�I���g�ׅ��*�@�_äg�I��`D��k'OZT	�@�t�rSaSX�;ė�<@���$g�"����C?~�5&��ڣ��V<%��e+��̳.��P#xY��F��(�_�˰�uBFi��j6B�?�6��'�?@
�����91���Q?(_��x^�S�I��:��b%_����;�6Xٲ_I�z�֢���~�w7�����r���~��5�K����}$*$��>�D�ǽ6z&7� ݙ���(e�~�b�M�)�����?��Xi��-��R����	�ݱ�5K5��*=�~��DdCV����1�9�a�f_�[
���4醗}΋d������h��,�Ơ5�"鍻'��X��������.�DG'R["�aҰ]���P�JF�^�Z�׆�З6��5�jrW`%�#h͒m2w6;��+0��<�	Ѵ�k��|�<9>��H#�hi�ٻ�@�{9e#���z��%T�����4K"��hn6���#���t�� ���ӓz!qPNy>z�'Ⴤ�VR�}6�!s����j,;�Xa�wZ2"eqH�R�SJ���Go�	}͉n�������))h{����k2���Ȱ��.{�'�峨��j����C�ى�r�o.G\��I�8��,�^���	I�o�?>e��ڹ_g�}3�ew�����p}=��i�w=�XJA}�iK���=!]�
��6TO����e��e���p_�yz��?���p��� l�m��N��|ο%���3��U�����Z�n3F/�Qy٫�.a��Uki=�+Ccp����	�*D���	T���R����	�I�F>[��OF�����:S� �#	IRj~��f�Hn���UAm�G�r֜�clT��Ɣ���7U$�sא�l���ܾ�r�Sk�$���� ���M;`�N����J���%�w!H��'}��(-��L �f�yG���}UTR��Y��r�h�������C]��V��)bA��
Ηy��Do��(�a5:�_牤Ə�|����L{�c�z���h B��Jv`�E��Õwv�(O8!��6��S�>���0�F��T�P%�w����>�TH���.��*_�����}�����fZ��Y몬۴i=��y�$�-����� e%%W�{/��Mw�N�������������$����6��K��"��%�U�TD[�M�~_�QIΫ�(,��m�冱����T*���ŵBq�A+�%ǑZ�g�sF�v��"������h�_�X@(���[�vj�|y���uH'}��E��{-�zv��]�q� �������_ח�4گ,�1�����@�{v��K���D ���/�Y����A������x�l�oF�����3lE1G"�t��C���%�/�k�Õ] Xכ�'p��?�忤����/|�yڃ.�8�lĨ6��).�#!�p)&-�`<�cS�&h��r�*�3m�ʵ������D��WD�1:��`����[[�̟=��-��Q�)�p�����Kbrq�!F��>�m��(>|?!%'��B��(��b����>7v$�B�3Yu�����Ž�ǘ��F�n�U�Q:Z�{��fM���6���W�y�0���u���{���ұ#�������{��w��B�Irj���Ht�Q,]�x��AE��9����?d̈́�h��s�@S$\i���P����C�g�Y���K��~�=;-y��u1��^�~{
�2D@���4{\�|��x��Nl���3�u�:Z������"M�h������̷Qև8V���C�ҥ�3�����N8�{�L��2�G���*p}#��S��|cmٕ�oS`O�1��Q��l�6�R��A,-�
�:��{����+'�!��~�3�4�W��/bf�*( ��Ջ���$��V��[O�i��Z<b�*B���r��6�᥆�+��7Û,I�cbb�oI��߈l� ����g��m'^FO���oty����ˍ5i�s��$7�3��JFX�l!�쪹&�A-��-�p_��:�y�d��hE/�V�f��VCx�����2����4	ȫKƸ�9aUD�U�mRi;|��Iji��}���o�XaoINq����'t�*�	!��I���	2��Y(��U�w�3^��=n��y���;�X�GW��i�?��֦�B��z�J�>��9@z�~�y�����׿���s��N%8TZpLhrS�n�7ם~��7w^�Jbnf+��f��f��˥5���"�qk���"md�(�VKeнф5/ԗ:?���G��M H�\׷�O{�B��o'6v�ǢCVZō1�#�.�O<l�8�9������
�'���wD�O�T����m�G������#�XD��m/���垆�Ӎ�����Ƞ�~d�	!�^��}>D��K����m�Qq�1�Į��K�6���AD�Y��}��'v�m�'˝�/SE��M�Hi��S���!���{'{�L��7��r/����r��7���׫����#�	��0s%jD�O'��1\)�Vfj��&��9� ?�o�/�wS�c����g&B_����&�;J�^������|
���G����ή�>XS����g.��2���|�GJH/�e��CJY#ğ3&y���Y�IzR�������1�ػ#���E-���a6#�,�拾�0zU�0�� 3���X~��s��O�2�I�� �!�O�|n@̢�����Ɂ��?�=�����r�p���+��H�U؂�-&��!l�.�j	�o��H��~cƟ1�'�i2�-T&d4�4ӷ�Ѥ�R���ƭ=��������]��E@X��2Fn�V���VІ������i�Vv\�x)n�ζ���g}`���p��{�bחʶ������HA�35~�E���dD�]��R�#� .��aa&���Ɠ$��!�c�h]*"��EJ�[Z���ׄ�lK�57�݊3�Ņ_�hDXPII���{U7>=�ou��/�+�LLVjӉhԬE>�����R��x��\>,Ҭݨ���A7�����E����8̛�Re��1��\~�W�U�\�a�
��^o�ri(p�_ř(jݜ��/~]4>��;�BS�z���(�I���W��S=Z'�r�kQd�uhE�l�M��j��>�Q�&|�_����l��,�s����"��v/8�no��I�E�W[�]�Mq�˄*0���v��v���eһ�}K!�we��Q�I3�E�1�W��%D���/5S<���k�o�H��#zi�(�Jʎ.��u�'�W�/@�6�jq!-93����������G��Gn��D̘�6rE*Wtj#5�`d�OE���P�/�� �����	U(��BRv���Ф<�+�e$	w}϶�IUGHSO�K �ʐo &�Fal�0��{��d1n���/}����C�#3j�3B�q�Y�"�YhP���4p��ګ5���D�c`�훏T��eچ&k�]礜��wa!���^���4�+E]kj_�M�.$�8�☊j��ybm��4e�e��o�����c_v/|5�)��M5����~�]A�����M��r���}�M�ܹ�eA�>���Y�MB�{��!�8����sh�˕u��2�<I�/%W��P�^�:d�#� s�H�,8����)@��g���r�q����c��
-�A8?�#��5(�O�U~4B��p�i/�-�C��焤;�5o7Y(.��eXc�1vޟ��x��Pa��'��4��%�y�0��Q�����bFkS{����i�2Ϫ+˦��Ĩp�g ��])�t[���!������H�)��� Ԁ�yI��N���ǒ�Ui���u8R�X�����n}���S�DŤ�L3�f5��wX8��_{~�G'�0�s)��|�% b(PoJW1Fj�_8��=�d���0�Iu���ݚ�H��)��Ϝ��wP,76�]�?n��N^,<"#Q�7�4����+�岅J,j��nl����U&����$�=a��\%%)>�'�d�KG�{S��$���ʌ*�$[M_W��[0f�T��WC�P'�!]g��mi"����[H�~7b�0�����5q���}C�7s=�Ֆ�ڟy�Dն��]#�"3�""��p�7��b%
G�l���RM�6���{���Y�O�=>��u�9�+�1�����aAQfJ��aJ�����_ ZEF�ד��.!��K���/��r��O����U.�NqI��6�;�t;�땻��%c�0��>̝�2�2<Cݨ�G1���јS��C�<5�E�(Ig���;f�JLW��[4�+����#=�p�j^tۊ3�� ��D����/��`	v�W����;�Ş��x0)��4/��B�\�.�4��_�&@�-�p	�ػd4���m��u�C���5Dz��tŔ?T��g�[J���Z����[*��ؾkM+.}���_���$��[̆m�|~�H�(�B��{Thvx/��IQ�r�~��[[��-q��n:�$�N�Q7���6�� i�3�#��fȜD�S<��Νy)�:�<&��M���s���zgtV�V�2������U3G��cJ}�������b�fiB.�w�����_5��O�`* �!D��j%�4��1$�3��0#ѝ������*os���e�;��a$��6AԊ�:��w�bB�W��zlj����0tF�4�J��(V~k��-��T�_�]�'�ͦ��G�-OfIeDT���\L��k[)�����^~��.g>L��Q�ةaˌ�g)M6����\%dnH�9В��e�I���G!��	��(� ���Ou�{���l_��Z�_�S!C@��u����:�Ϲ>�r�
��-���O*)��.�ֽIO�i�p�q�$��˾���,�XsZx�Г"L|E�������à��y7��'o*�5s�Sf�V/�Fy�9q�t3��?��	�%�?}	�=�����z �����������gR᫅��eq���͍|/VĠy�:�3/ �cz>P��_�p_v-�L����|��o����Y6,-��&j�8+ve��B�i��#q�@�i��]?{ �a�[���e~E �u�(RW9I�Wʤa.�Ĉ�:O1�li$��&��(a���J�����ٖ�	m\�$��<$@f	Οm[&�;b�换j����B�/���ET����z��pB�|Y��� ���X�l��k����'��[�H�ou�>�,�ON���'�8,[֐��Dg�V6D4h����V�1�\K��q��g'坮����W��'�|\����|X�	o���j6V0ii��Bk�������Mc:�z�%jKm���2U�tt�%����3��[up7~����(�Т!�QY3Z@�S<C���;��.�\�s+ծ"��[�)m�:V͛#|˕Z�ˈ�D�@>a���n<���੧jv���-���O6nS+�#ф�׽ ���?���g�0��,|�.nc0V�)�~(��t�P����vpk:)��tIԞ;��C���yK��$�bI�%�������)����5���-"���g����9�`���v1}��'Sڅ�`�ؽAW���� �z?�.����o�� Q2<y��
���$��'QI�ŒL��w/�7�^���GsD=
-��p��o�3��>W��J�#�^5�s��A(��@PȆ�P���F}�ˏ��l%��v#����a� ��R �$����}�2��ccn�=��82����^mu��p(�w)Z\�;��ww+���Nq����;��������Z7Y'�I�ܙ={�3�K)A}N���?1��h)D���x��Ev��a�0��X3lΟ=߀�[�����Â6Zr%Ybv|�=v."os;6ːs��8.B�3~b،cT��n�τL6�H#�e�[���'«q#�|�NkSA�XE6��zl%=���b!3h"\C��{6�'�z�In$Z�%����zt�;��t��o߽8��y��*��䞷*!�X�ٱ�*�Koż'�����b���)�P�
ee!=[�1�8��-����z{{C(�^����M����ި�~��\�br�j�t�sN�-I��`�����e��x��ȓ/����OT9�z@D?w��|9f�}���km��p���L�,-����	��Q���]�N({�*^�����Ći��9l���v�P���6�n��m��Mz	�N���H�镅���#�-GV����
ѻ��1	����[�0V�� ͷ�]<�y�0S5���ɂ���?��0Lo�ݿ���,'�#��v�Z�������[��Yb���<�%gZ:��H9�bl0{k���K����j�iS�+��E1v�����]�q����L/Z9����4(�}���!O]�|��o�}�'�� jgԆO7�)Xک�l��i�?*{��9�6x���
��E�Ĺi!�r�-��??�nsB�.7�&�M�D�Fl2P>�p8��j;�V�Y�.YBkJp��.E�]���	ҏ�Ԡ�G�hUqGk�\yt�s�-�>v0f	�B��֖��ꆸy�u�.�r�,
;��:�$�}>F.��@� �c2Tc��S��Ni)9A���H��z_o(�:= r�|P؛?λ�jLpi�t�y�^NT���n7�T���M�K�e���M-�>P��9+6�P�?g���K��g'C��ٺ�F���o�$>2;r"W��W�k��	��݈`���`�L�y	�P�j?��T�9v�k�֏-\<�"��ڨ=L3_���y���[�!��SG${�"�ɯJ����v�#^5]��5���&D�U<����i�r;V`�s�
��{G���
����0����ބ��L�g����|�2Q�v�����}��_�炃=l��>Gw@��X᏶�C�{�݋p#��m��;fy0�>יw�&O\Rj:=�0ȷ�u�~ϱ��3�4�̕+{�t9�i'��)d�v�P���V���*��ظ�̔T������D�eP��F#7�]�>���Ǎ�Dԡ�ғӁ͘�����'}��2�r�2LG����j����1i�V�?"ѫ ���g^+��{3S�x�M:�S�ܡ�c���n�Nݖuۏ�(*cy�+:9h��{�d:��Yh�@�Z�f�Ew�$�^L�tԜ]�XX0h]���SL`mOB��Cr*#�hbӏ�-�w۾���nQ^�f���J�{1>+8��T��ZZ� ��Xs��c�{f����X��7�9U�cC����Z��Z��4�URq��eS!]4Z�y�eC|��R��� `�%�Ƹl��^Qg�m9����T��	&<�&��[�o��`���DfL�;MK>��n���g������V�bv�y������P;S�]�jED�p�z�&7�_X�6P�1�;U"4�[&-G���Ӯ㺰scN��{�YV�Hj�FP�;�+76��kw~C�^�ɍ�V3��p^� ͕3�?����i�O-���Wh]F~��[�@�<��^�zG3?����Z0#Fn�ܮE��<EJ�V2�bs<Q.���rV��f3�"�L���h��1C��)�oo�{�3:A-��z|��JutR�cpd9��7T������]�ϫČp[�`�Z�_޴�;��x�wϯ�=�WV��r��L�1t�Rg��3��	xd����^�\�E�CH"K�z��=Ҋ�DHI�����d3>Xә�PѨμ�yf�_�16~#F=V��/P��0�Y��Rjؑ��d�ӳm���y��ˤ����O��C��O�O�c%�3�o��iz�k/r؈x��%���SY��v��̔=��K���o���O8j�FN���fi�Rᩂ!6x�R�us��\��l����w�\d�4����UT[׭3s~҇n�ŗ\|�?�E�,9w��/�C��h.�����A����e�fb���$F��֌_�Ɋ�|41�+%�����::o	�K�����jB��_&)j@m�e�v\���x��_�@������0�y���g �J�b�lٙ�Qb��e|�bTО5���J�H�g������0�x�w�D��<?m�N�yЉ��ӄ0l����F�����1��5���=�@u'a��(.�*�x�6���_)q��͛�J��j���[���4pbBZ�����G� ���d���f�v���dN��\}�("b����Dq�4�`��7C)2H��Pغ�����'ע�ƕm�\�c�;p�%*S���?�:އ���ο�ij�㘈�������Dӻ�����`�Av^U�����y�Q�3���"P�k9�^vG��@37���E � |ئ��v<J�e!�F\�W�2  ���	P���h�U�u\]�v,d� 9����j�3�|����6��/w݆GK�������R���3�#(|W�6l�]�#Dm�C����L.&��>�q*�?� 't�}VRB1v�oɓQrѻ��>cyz�.�v�^Ptu2�F����~�����h�G����~�����L�^M��F���F)��8�? ����ظ�災#,��A|<П(���PV1@Jf����? ��@���ʘ�?���%6��]��48�������0���$�I9��)����vﲇ<Nd�C@�0`6��$&��y�[FQ�f�����c%;���ֈ���@�Q��a�=2O�k����%��N��OҠ�~f��%`U����w�i�_����{+�j嬎������܊CC"��'62�\Lv
�iSF�U<4q,}�?��'��B�`�Զ�ZO�/'?�@���j����hh�v��rh2<���N�e�z0ꓒ�nTn��s��~��G�t(k4��)S�R]����t?q<���o#U�b1I}u���u2��87��8`��1���S����+�,zv��`SZ�5����2��c	��B/d`4
��퐷�/^�H�0
�7��[�k��,Ab�`&��C�с�i	�=}$��n^���d�~��B��������*�����^���	4P�fI�D��}B����"j�Q�,�1�5�"b3�,���Ql��/P\4D"7ȼ��OT�������uǄ���I:�-���X.4t��L�7�*�g�j�Cq��f`A���(���@����*]+�����D2�O� ��$�a�ָ�R��@�"��#P���b�d� ��I�:�ݮG��ɱ��\;�ܹ�\_/��V��x�6ٕ��1Y�x�?��g�֜%BtF,�g"u��_�8g��q�(j��u��Qjd��-u���6��Z�R�#Ip!��(jE�ǃE
S��p�E�m�vb�\E�!� E6L.�����`��_�4���d��E/�Q��.�,�H�4�n��!&�|Swsc�yV����֎��k�&t��hi1dT(<;$zL���j�ͧoa���]��Mg==�����~V�M�W��"/�m��
V9��1�	w���4��9EP��C���ÑaC������k���a���%b���Z�
����������,�!��EaJ�_+���7?Z�{�S,>�}�^a�k�80��ml����O#�b�⿏��p���JI���o�@H�YHrr�_[��J�	#�����$�=�޿�)���>���gP�tЂ)N�����͟����l�������Et���� bӵ�mp$T9��{��)U�X�ʮ�`��g;�L�VA�Ҫ�Z�!	�Ղr���V����`1:�p"!n�
O1�aYmu&��f|HW)	2�d67��V�]`�U�Q�A��ڊG3!! ,Z���V���G��Ǯ�'j�����m�ڑ/=9;/���V���R�瞯8\Wk�P���>\.1k��Ng��f��a_W�J𳮢�p��Б�	���`��/Ɍ�\�&X�L(fA���%�����WNc&H�tC���i��!2���Z��r�Z��Y��=�l��.�\�+��-��$ґ��6�_��������b�R�;ʾ�^'������*b�#~��9��`����g}���V���HF9.d�����4}��[mgqtt�Q��?�9��ɼ/(赵����j���.��ʌ_�mİrZI�4�>��;����<_���@E[n�ڶc�m�
ϳ�f`��p�F��~�3[]�=m��[�d�"1c�;�t��l�����c0���������^����/Om;%]LC�j,�)O�����z����Ԣ�#m+�<}n�]e�ބLr@��Pf?��l�U|�<��1����P7�}c)��O���C�5ttI�na	�.����Yr3et5i9�o����'=:Nb�����s�3���'0��^F�^D�J&�E�{��K�6���[�OV�\�������P�Hez!��*Q��'�\���P_k����ls�o/Pb��͎j9�E�S��w�Ck���=����٣�C �iy��f	`�pP�p4FJ����lU�������7�g�r��L?��2g���������p��*)��R�)fAV��8��Fm���ݍę�t�ޚ���!�'rc��8�y�k��Yw`o�[8LC�)N�[���� �.j�]h��)�\���'p?�`��A����B�%y$�����g�����cT3ɒ��*��d�Òk�ˍ�1U��xl^�b��"M�r�Z���z)S];�$���}|��1�%��GY�XE*TH�I�I�z��N�w��I,y<�6�c�j��W�b� �*�x!�C0ʦ<��$�f�3�������z�xVC!��rЈ��0����$�;��͛$�50�ǋ6u	6��"K�l�梍 Z��f�^hF���\�{�݇���J�
W$�p�Fܿ�j�3�9�O�v
<h��5;�^l6�jG=�#�đ����~F�R�]�
���?�͓�(��w�yL(NY��{H�b0l�2�!�!��
Ж�]YAr�ǒ��(vG�s����}'���/Ex}�r�HTU���q^�{��[�"c���'�?P��;f�/�SY�_�����лv�t`�j�4ج9����+U%�,vȀwrd��Z
�~���h�H�>e+�� 7�t�h$�.!73�}����ľ�"��q�xí#1]�������Y���u�������۴j�C�!�~�������屇���r!�9�7YV2��p�M�T��/�"��yն��8�Efn�>E���2�1n��� �9Z��?��v��U������?�Yv����Ax��G�x?��.�6g�21,�bi�e�N��B��T��:٬���R%F*���9˝՘�G�d'A��dH,���dS�c�)�N��N�Jݮ�����B��?���6S�6R1�"t#I*u�<�a;5�,=�h��Ѝ���
>!u�z�Hȣ�2T��ڊ�p����]�\�}��\*���jSܴ��� բ��Jv�54�(��ڔ3�Z{03���8��	�~���#���N��V_��r�ӂv�� (@=�������n�{�a�|�$��t"8c��3"Dָ�-{8*��u�<�/2�(B0d	z+�y��Cn11��9�G���uؤ�f�Mˊq󐺀���о��L>�#u~g�5��'����m���:4��G��m0Y��k�_�_���<O���j��ck:� �9�fΝ ����]�!���0�~�l��u��m�&�
'F		hT���?=l�J�O	4p1D5�g�^�M,��m����łK9(����G�*X�!r���Z�zަ�c3X� px�� M���������G6���t�~/�Ux�빗�D�õ_<��c���}��*�f���o�����V�!d�:k���#=��b���⬽d��}qwG�?��q���z�=7�\s���pa>���yic��2���}o��k]����<M���E^G�$���l$_hp�?�äa!�x������`�M�,hm�=�G?\�	���|3{��A���i�#�0î�����q��Q)R1��HG�	F�g�k�]�oÚkٳ!J�F|LF2��l�Y����f���K�)?��v��	M�1V�;��7��XhYo�mP=�i�۬=hXC���$`
�(���	��~.0e�2S1h������";�Q_-�	�4T��}��b�\[$R0��H)�.kB��V�j�3�jeU�b��T�ɍ;��Pg�4mC�"�_��x=o��:k�"D(ɶ,/���Zѕ8JY�4W��\���� �6�����y��v*�����L�
 �r�k�������?�:Q�mL��w�R���HH�\��K�]��1o5&%[����D���~&V�������h�f��΃�i�йSn˄��g����}�e6�Y���ˁ����l���k��0�q�d�ď�:ÿ�t<Xz`螏�i���U'K�~�����ss���R�Q0�,�8�d�FҦ�����gw�Z}��Ai�٢SkQy6`��̻�8�ٻ&E$ɱ�[�q�V�!��q�� 4\�f�v+�@]���_�*�;��b��&�3I�rw�^8%��r*{��it9�o��0�����-m[M���w;�?g�Kψ���6B��BUZ��bd�	H��yc�s��*�?�.�}.�_^bT!��
�2���:^��s�Bl�r�� ¢>�\f�]�k���,���Y�&E5r�"������1��b��b��P���z\=�ծ>鳸�X���Uh]��f� ��qxx�b D�i�%�elDA�[��!�����!��i�|¤e�s�4f��XD\<^:	چL�B7�bd��֦m(H��ܙ���n�v����������vi��o��Pa/b�'�zI�s�B'w~.���t�o�,)/M!>���pIUS�יnv/3O�S4x��$����	I�ts��g�;o99]�*����۩��uIOCH��m�o�8rW3��-/N��D�L�~7��������l|S�ũ
s��]�7L���! � k���� ֵ����ID I���g�Q9�P��˿7X�;`�;G�{���O3�L�_��џ5��%���P=�[�rq�;��l�<OĜ�t!�Ћf��ٲ�S=�|5��qcA�Z`�KXD:í�1F0>T%���4똯�6�8�7��P�2M�����.FT�y|�����`3A�]M��KpX6b�6tC���u�dH���;K��9��������(x���M�����B"x=��I�Pl�;p��\ �L~�X���^�KΘŭ�%]��1g=�緍4r��rjѝ���g��9����E�GZ햁���L�� Ka!��Z��p:��ߍb)��������DG8���fg:˦"�>7��k���r�P���K	8f��{8\�^S���f�W�,�x�K˭P���H	�@5��9[q�]��%"��E�'w�V�X�o��D[w�nҨ��h�ݹ�LdzC�����Oj��|;�X���A�c��Dm�e�[�|�j�$�TCE�4�� �c�&�f�L�@��i]^G�{�C
�뿸�W<_J�#�dK�g�5/g��/b�&���VP* yC��;�l�HA`��S@1=�ՆL�e�gc7��v>��`{N[�a����jX��M�{�+�2�8�dg���-Q���)_�����W�zb�e��,�����:�r^�5���;�
C�?��ϰ$���4eQ'K���c�_�*��K�	�G!
�����ô��P	g�S�j������
�A���5E��B��;�L�7fH>1��؍�%O����˰���zSPg���&���ET/���p��E#�u�N����Q�&&P�I��)�O1^����V|䳡�e��muq�Уq��R�0��ʰ��+��ҥ�)`�]Ğj�bO���f�6�N~�f�u�`��ui�w�A�����A��m�6�CH@R:O|��_�Kk(M�k�ά�zRv!��pd��~`�~Sj�'C���Mq��Yj|�<��	��5��9 �m^Q\�LbwvGm�}m"�,_V�`��~�9�����rA���P���Y!HqM�L�.��b�g�j�P�:��L���NsV���:�R�}�Ψ�fe~n_����X��̣�z2����@s���	��k�N+��y�����M*(Z���tN��m�?��y�~1fd0H�^���^�Ikm9��1�=���1��g]��%��j�-�SY���ę0��,{��1W�3�C��
|E��s`����9=��~5��&����T��)�����v�L�r8�MB
�U��#�~���."�.��2��4����G�><�A'��p�����DC+R6�$p� i�~).���Y�'K��H�'V��v: �>�����u��@pr�.�T����&�Ўg�nA�qs}���u�,2��q�1it
Պ�ȥ�2�/jcq��hy�$~��9���@�G�J���K�������e��a��	8J!s���n����H�4���q���N��֑Y���y ����W�z	��n�W�l�������L���|GFU��{(�:P�I�]I�+z���c9�^�;h����|k*fx���6��r�0��Qb���B�;s>��������t��C�lE�P����UIZʣ^����#G���C�g��e���:��vb��a&��7�o�"�G�,,c��;���T0OZ������G[���۸�x�}Ӡ��g'TCD#D8�����9�l��/7�+�,'൚�Cy�r}xpi|e+I�_���MC��v�X<3cH*�;XA^̎�j���gr��D����s��L�鄗��D���k���C��~�97�qbN�W?DĒS67��5�w� ��0�uy!4T�/��b���� ����'kw"ˮw�����g�KF�.�E:áԹ�|��R����y0�T�ώ��4{y܁��zk�8<��󚸑�;"�}�a��U7ΜDLmD�]֟� b6�"'�W�+i�t���:��V�w��V���f��q�S���׺�O�"��6��;���:go�,���V�+��t#��~*����?���\�<n*MkE�	�{�k��d����vޗ׫���˵���q�@�W~Hu��1��)�hrR��VV �:3�e���Z�j�lvŧ�s��#�%o���U��}���S����+�N���Kt�)�?z�0��?�M��v�j���_���y~$����o�߂�}W�~�Q���N强�� �cy!��u�"m6�:�ԟ������`�4*2mD��3+��lo�qa�f��~��(�[��/k{��|a�R��y�c��"�
�rCw밫��Rh�d-�Ѧ����ve�h���~sb�l6�/�#,foÓ���<x���36��+��V��l���ҦbY�*�Z�>�R��!~MC����g�ԙ�uC5;V5h���𨿛���4u�ӽĄxLC?��4����g���c�rn��5����ݬ�]�7Ý!.��(J���T�vD�#�8�2�ݢW�,W�H!�|X��]�x?I).��������m����ڞ����J\�@;�_cT_��C��F��k��T�Bi��_	��wMX?�h�9��݁0)@��{�<vj?k�!|�4�IM��!�hȏ$�tB'�u�+X;
�(ӽ�����]��ܷ;!�2�l���6B�MO�L�P�ʬ�}�V9��g��r~:�S��PN��z��9m$�L��u���W��"V�D�w�:�����T���
�Bk/�L�ґ�ty�=�D�rBa�'��N��Z�j����J�C�d�?jH֜e{8Rv/�'V�U�A
�O{F��e�;Ĕyx>>x@!��ʁ��|Q�hO�� $F䟓
��]�t���IE�f�:�F���hr*�,qʑ{)O~�9�#O"z	X��Z��*�`݋Ta7�z+�͗��g{��җ�؋��КV!-��ҁp's��|���������C%Ae��wA�=�Bo:�z�Ɲ�}��K���b��^T�4���ٻzں��w�P6V���\��]�ñx)���;<blȵ><��<I�J���5-9;F��BC��o��:��7�uD�ۃ��x�D�5[�}�O�8�͗�E:v���\����a��3H;�|�rwU����-����C��M�Q�tKa���XM"��I���1�Wk�$Cۗ;��v�w56H˛yjۇn�}s8�Ϗ0����v����fw��z�N�zh�� 	X��x�M����*�̓�+T���(\c9w4�u/���dˏ0�P��'��p໌-���Fo�"���J��ց�s�A�s��}� ��-{��� b?���|�m "�1�A�}���U[ ��@�J�s�t���@�����3�Ƣ�D�B���r�2��l�P�"����6�2�p�'(�� -�rYK��r�y�ԑ&��j*ܕ6�Wo�]��6�@�����"c����óEp���>ވ��_�����9�X�4?�äg�GAA졁��&��jQ?$��1�D����ו�9�]؇�WN�I0�{{,d�ؘ�/�x���V���ը��7w?`Q|�@�m<�p�,�nOX�%�s=��b�"�aY����B�KO\%q ��oqU>��+����d���X������Z�v�H`�-��):�3����,Z�Er�r�$);]Rn���4��3�������u�tF�uwJ+�i�q�mD�jܯ��_�����NQ��&.C��h����p���O��%����˵��U�E2���VOs������}���N�2d3�����A����/|�.��y����N|;�+�ȳ�Z��!R���/��E����JaN����x�fg&��cK����ܛ<��.��tƪ=ļ������S�M�b��Qs>X�|��T�`a�_��k���7�����1X�����{)�1����h0#���f#�����]>���L��Ͳ��(����^w���7Oy�~�Fd�i����x/-� 6�8e``R�#<��-{ܡC}j����E8�  QX�+% u4��徵��� Ş��Fy�ss���8��q�����^YO d�Ӂ6WQ�xP�.�]~A�v��N;.
��~�m�y�iک|�v�rE�L$�Uv8B.�� Jn*�c�g��V��<�	o���%כ��wOȏbh�ǹ�F.jc�ݻ���;V��g�;�������]�_�J����GF���c�g[H��D��M��";I:1]7Mu�L�s� $bFZv[�����+`��d(������;-�S�"��@�I�QƖG�#ʋ1J�`!�T��Ґ�˒�-�˓@u���$��L���7�E��iU�f������*=�e޽_���Ȼ�\��@!���I6b�2���f5�8G�� 'I�p�1i��C�%Ռ��s�������v"��,և�D?�D�R��;��a�$��@��� 8�/���T�c'9w
����p1K(��j�ʅC�"�M�j��o��i����s���m%A���1�Q)��9��$���L]��dX��3)�������4t�BO?���[M��я�����S��m�;c��!-�MH\S�&��`�φ1���7���jh�o���Y�˹����G��<����^W$�AQ������S-zF���.�w�ԖG�a������,Lc�4��S2��gF3��WyT��J9��;���&T�6���� �c�`��;�03��k�����ړ��*��a�7�s�Į�|�wc��J�t}������ʈL�x5z1�_I�v�������SI�1+�o9�Jb�;*�l��T�9j�Z\wr�$9��v��u&��գ�t9�K	�;�; �c��`.�H���:L|� ��`:�Z��<���7hhRc��\�5�^�
���(Y����X�d ��>�����(|U�RD���ɬ\��)�ޗ���z�b��X��1C�p�B��x��ĭk(��<�����<63$��_��D2zTy
J]�[��^�)���ZUؖM�x1���#=�H	J��9�XD6���f͓!�s�m�#����a�G)�����14����o2��-{�i�acVc��}��	��X��Ea�a
��&�XNR=#S�o�[>�*��amxg��//���^>8D��~5µ.G��1u���t�����j�hj��#���M�X�[꛱HFnn0g���P�:�a��0��7z���X!݁-?��%���'ȷ�|,p�+��lhz��8�+̥���oP7�=[���+_F�2����8l��l4�Ud�ٓ��~�-�1������aq4oq�!oEm���_���I�(�/1��⨛�0�	�G�7���Dv4N��YL(�v�9��4!_�� ������`y4�/%c���r͇hR
��pDT찪)��k�e����4���>M�#��`v���0fh�Z�&��l�)�0��qp2A��X�#��u�k:/��Ze�Sa�9��;�m��������~�>�杋����p�$(HsX=Ey�����%�@C�
b���̖_[�B[7����'>(}0J�t���l���0̄�"�й�6D䩔m�F�j4Β��HvuZ������I+�4�7�^]��A�'##5�7O�M�T]_�d3��6����#8�h�Lou�NE(O��Ɨ�0M���3W�S�,��C#=C}5�ȇg�8��R��9�rC?���KE�V���2����w.�>3�g���#�X�E~jnJ��r�|��.e����b��n��_4�<Y%��۵���\a:�e����؎��_�M�Ϟ#��o,���G�z�(�� r���	��
������?���
,���@VZX~[����T��=�;�kl5^A����.�0����vR���z��:���,�Hx����']̜�oyK/e6�	Ke(�:҃#�i�ҲZr&�d52Y�7%����[ǽ�N��_�-H���!OH�����x����C=4
^�\��UN��q\Q�9�9�iJqG
�M�_s�=�>�^���_�z(n���d=\�0���1�Q8�쀢�f�A(�aLU��,L���<H��ۖ@�+��P��J��� >��BAr�VhL���Q$BCk��c���XD���yA}�î���oݥ����i 1	�����`p��/W�LH�a�vϟ`�}UoS�4N�-�å�>���W�ݴ���H�B�=���"�Zr��G���y�&+��q����m�GylG=����%J,����fG�v����>�&O�_X�D̈́�eS��8]/���0�tSk4u^-`���&	�\G��Fہ:�b򨡘@�>8P����g��"4'��U4Q�AO�CR1���>I�|�_T�w����Km�*3��GI6�0\՗�Un�����ٔhՎi���y|?]ws�6K�|���k?.]�g��0rع	���'����z��osq��bl!��������_P��K�r���s�x�N�o�r�݂I��N�<l��S.�fΣ�܅�S�knWI��op���&�A��{ԁo����s��#=;%�:���C�<��6�h�b+}�Jz���
Kо�Z�V`��10���>�w����
;���$�s+�:����i|G&�W��V��D��}?-;!FW0m�|SC���Y|�Y�n���8"���f7��/'�^� ���ص�P�mnME�}P��XWK����\�ʄ�oj(EUc����m83��m��ah�m�������@�`(K��L�L���x{��e{�b�ך(|�p�N���͈ɧ�B��~ȴ7���oS�s��{œ�̳�$YO]5��Ŗ-�[�Z�q�d��;���(�}���|^�@��q�A���@w6�9����#Ux@� ������������g����Y۲�̸���:c�UM��²yy����(�~հ�����e�^����
���èp�KLqk�n��j��w+�1������c��˅v�S�Skm�B�)�Ђ�#qf��i�55�ѵ�����&Y���U&�z|�7g�4��H�#�!}}<.S��v�h]��Hǖ���Wb]]� ��p��I�g�F�n�Gž\�oT�!�+�g��܍"_�%����2��țF�_,�1Gr�<�}��xk�X�K���~�r(�d�	�{Y�ho��G|fN���Z)�Ǧ�#de9�\��	;>���f`S����EL��U?�S��B�7��e��p��~w������SU,C�_�]v���jw�!��D���m�9X��i�@H�WH��~�����m|ʍd�~s�#������כN��><"/ �m�'��D�$���\� �?G��̙es5;�b�~3���|}���Q�l~'o��|�����08*)�Y�%��@�߷9��{ŉ�%V��ƴ��4����i%��;�y�N/���:�8.^����Q���f8�� 4d9���I����.{��5����
\v�y�������,M@�=]��f���hy�ԦպF5�����;����uH����I���:bQQ�9N�����ß��|�Zo����հ��k��וu>���ǟ�h%d]ٌ��5��v�	�u�i`�oU���|8�,���v��|ђ��\�4�LUA ��1z�r���!�g�Q�I�6��I<]�����[�.�9ʪ[�����M�f�yÕ��q"�Q(2�F�	�����˻2���·���+��bv�|���X�o��a&����x��k,g��d,#�K21��A,���w�Y�J�l�PP������JHj��-f�q���0?�6i�'Q0���
�%e���Y��f�~��w�c���;�!e��3@l$�r��׊H�ټ;�x8��(��6����Q���Z�Sl��X���ؑ���;�����!��Tj��]c[���4�+�ޒ��d��b�Kz^�ļ�=^�#���qh��n�Cm��c�r�E3�<s^�9&^	R���UKo(�1�D	�����z�b�dI�$��j�����>��E��@�"�4س��r�X��5˺�N���3��b�����n�v�1#c�^x����r��
�T�����OP_>^Y���T?M�EAt��{F���֧(�~�+�� ��Lp�V�!
)�t��/[Yo������(G��8O�1��Vd�1���	4��! ��w�tz�t��cqB��5�aZ*�jU drBi8JZ*<�f�QԮ���;{0zSQ�1q_�%S6��ׂ!'����ȥ�P�q��۾֡���?E�i_��x�Y3����e��u�_.�>�(B��D�&�X�Aj/��$������TTĊ�|�EM�W����/	��,%�'Y�T��?�i%�P�}C-�y�8��[ֵNW�+d����٤�#Y,ꑭ>���2Fd2c��YݟF|����L:*.��b ��3 ��i!��S0�!��'y�Y�*!�ɑ$Pk����,�]��������|�T���? J��NH��E�5��E��.�>��Ɓ����l�a��Oh�a ��ȕ]�ќ��>M� J#}dÁ�T�00XE&@'��L�V�X ��P������X���d��:�O$�4��&�0@|����r����x'u�ǿc�dM�yZ6�z���fZ1�CI@�R��=I-T#*�$3>��
�9(a!��	uZr	�ʨ˱Fd!� <=DQL���c��>/�Ke<�)�X��-�_9�Mit�a�PkSjjLh�)r�K�uW��
F��R�[��9�G�ɝ_ğp�)(����\������Nw"�����Qfrg��7d�y��:�S�nt�� �=�V�<]���b��x��2�-�)��Zp^��J)�D��<�8UT����H�+�p�"JC>�Uy���A�,���b��PX�f�D���:�h��ݎ%�S���eG��jUQ�5KŎ�KV� ��gv3�K>T1E4g��ZF�磙~gME��h�$&n",����֤�7��ݙ����3�yz?��'���g�)�X ���r��ꆪ���*.���琐L5��kƪ-��:l�b/%�l���#Ʒ�P�N�[�*ʏ��@��Z���h�-�x�)7� �"2����V�L��/P�~+7���a����i��Ԇ@�����4��JE��N�.��g�|r^��g��î[i��'J�s�<�p�~��*2O�F���~aΜ�g�Θt��@����jrs��j���F����8�,"� �?���-�&p�"444 `�B���\W�]�dB�=L����*È˔Ýd��!	G���)�����G�;8G��[�Nl�۞L�L<�m��$۶mۚض1�3�w��'�ԩT��;��׷����^)z�d7�Zt�M��K�7$8���\B��������WF�%N�DS� �W��gˉG��k�fz׷�#"��dz�d�`X�������wM�ݑ8C���v�6R��-�=Z�w�jڻC˄��!q��@҅2����5�a,e��f	���G�z�oˍ@��"�����#���Ju�A}�9>..�ޞ��'Z8A�Z��tx���G��<��d:[�/u+�nԉ=����Jiee�d�8x���_��$�P���0�mb�!y�9A!�/�S�t�
���
�^$M�r�a��00 B|�k177���H
�%nh*L�v���T��dtl����RmtrS!@X�б!�;" ȑ�bM�(.-M�׸'	��K�L�K}�Av0�$��G"'���UW���LA%��eg�{�`G��-�����u��BW������?�Ч�4xRcLW��w�[|cD����B��y�� ���a �T���D�A11�_�Ӑ`� BHJ&����,T�S����НVſGW�2����s�ϯ�0��:`�)��j���)��Z�Nz0(L0��7�熌."4���p?&�>�,���O�x@���O�C����as)I��7��Ȟ��`�K�qN],VM�!���N���DC۪ʈ��$(H{OJ|�+fۦ���o�����5����q�˙���W[wnM��It�Mny�r�U���AVS�"(�<+�ᜃ�t<�����]�xu��������锭���s�p�"nw�D@�nS��SL���i P�3��M%:p�\7TAE;��jR#���CRwx?-dp���Zz̏&0�4t��o�r6���}<O�j��
���7������}j�NM����'b �YDpz��eӝ�����#��I+���;Pv�'�e��󖢥�~���Dڵ��41M!+Ɋ�?���5�i>����J�@�1n�������s7�|A��O�A� �O�P�-�k]%r_�ȿ�}@�<��k�p�>����rk&�ҹ��ܸ=:愶y��9�QL�-�,���s�(a�J�#뽆2ಀS(?႔��9�"Y�h!5���$��E����h�y��6���H$�(P���s�2��y���Xn���c:�y&F}�)kJ+�r����-})۾�O�,��2I�JbP�\]��(j'�pJ�̂������e�P���w΁���,rU׭�rx���M�,��AO��$�
�X����A������z�;���8c�g��-w6�(��f2�+��עc�3ݞ<;2�J��c�����)�K�ժ^�S����|m4�y��	�������/jZ�%A�bnU��	nJ����Rڽ׺����ng�O��/-���o�N�]	�'���Jܓ�^M"MD���	�ь[E�I���<v`�o��f3ny�9���3/���Sc�BfM���1N���4����ު͇��{��5<=�5ng�;0��{��/ 8O��v���?r���r}�����AwȦ �)�����`���=�ʛ���'̝1��J;�������:yH�ߙ��r�s���,��؛��ճ�$�σ  ��'�_D��G��@TQ'\�ϊj5�V�8����?��e$R�7^2n񻽵�U����[3RK[cI������կ�<�.��������5�7g*{ktj*?��h6��S�#_���9�� ˡ��;��D��~�"��JW�G�����KR�Q�z��+E:[d��E������,��)��tٰ��ӏΆ�d�~�8Tf)��uxh��I�k�q��4֩?N�c6��^\Y�u��]$)���K@5d)m�X�C+#4�R��[`�T�����0���H��g�S�!����r�ѶORc�U�ժfG�RLm�����uآy��T���BqdP� 4b	Ԧ_1A�:��$9�燀��L�y�;o��[o�Ȱ_��r�a�^9	���NKq�&�0��$��NmT�����5=�����M��y��X���r�saJ�
k5yM%���d!��5���`�8Z�.3��ǄS���H�P��c1��݌H ��nM���0�ڽ_.����[��W VȞ5�?ʜ���/�#zp��"Ew��&�cE���'�PI��4����?6�n��
��a	�"Ǹ(���="���H�{-�C���B����)�YO�j�-��7$�B#�(Q,8HF8�D�F8�`��R��	υ� �#3���:�q5�$�j�ҽ��a��tx�n��{�<^���QJ�@kw�'X����p@�P�3=2Q�O(Ø�0$p����������Z.�6M;��k��o���#; ä�C�^�ls;K%d����x��l�y�-�Fu�
�寴-�T/k{G�U��«̅n�z��-��m���L&!�Hǭ!'(U��)bte�#��H`�g�	ոi�����N/��(H��grњ�A��X��"�B�� ry=j�I�互�}ۢ�?@k��u	QBw�[i�z�;?UDA��N��N�l�{~�9�k������:>Z�6��I��
���`p,��N�ǻ�+����rWv�1��O��(�������3Ո_�u�I0+M��~�+B������~�R�y=� a5<*t<��D#*�S���N�;�4^�����D���&'�3��rN'�B�m�@�v-��rPz���0�(r(w�Ǿ�E*��W���3&~�Ab�[i��V���ѿd�m��a�b�I�a�J�.�Pi�^������m� ��s�t6WC:�3�!�m^G��lx���.�J�[WO���0�ѥT`(�d�#�q�q|���R�� ﻞӾ�{B��z��f�q�yY�M'6'�«~!7�&��ϔ�tCȒm���k�E��ԕ��#�0Ps�W���bbx>�V=��=�n=����&Uz}���5�=tc壼�wC~}��Q�ߤ~7���>�4ːW�7W ��E� *������q6��)A��A*���]�RV��~�JA�C'�9ߞ���rșW��U;��*T�cԀ�b���Gĝǐ�����:�fWo�N�HK-y���MMd�q*�忞>���1����w�pq�[%̞���#�_�����2ZX�>\
�w�J�3O�����)F�ۡ�UT3���<��Rf����"p��RT�0�+Lǭ�3����od�P�i��Jwp��"ֻ�@��N79�ņ,e����~��)J������v�xY:�&�-AFP|��F0gR4��$�ȓP��?YL鸪��h��8���e-��7�h씵\&�j�:k�*>��l�T����C\���B#�F�!6ϩ0Jh>N3��6� �H��nO[��6Cڶ8�F�JL[>���;ο�h+�0D�g��`�����@^�3�͞s��**���_�h��=ϡ ��4M}�� �s���a��LE���DNZy/�A��+~t^*f�ʇ4��T��.�OˎY�������,��(�E�g[C���4i�hl.�M����5O�����I��8��PJEwx=�gz�k�@�UF}T��Y�Ш(�� ��r�U�bJ//~:M�^�*Uؓ>���r��FZD�}K����9wmT2RnK�Ȝǯ� �_�l����ƣ���/2.��!����
y�2�V\�m�	[�'{�� �v�*Zl�?�����oq�K�|S)YY�ۣ뛛�Ώg��؉"N�)\5�)���b��]��~�{��?6��\RbC����
2ѯܰr�������ch�U�b�+u��8>�ө�� ��e��y�7�k%���s���)
&�@gp�ٮf~ُ��׍��xf?�<���.$���O\���b���ܑ�����)����{�T���yhS���yݢ��[O�S�5"�<y����딁ɜ�.#��Va����֪��
f�`}\���#���	L_�hEhŵOZ:T�7n�'�F�]��S��ElO�B. ��JO8����8Ӻ��z�a�����Ew̓v��ِ��*�z���~Ҥ�޲!Ve(����q����.=2&���\�E)C��j~A�Wւ_u����N��g�W:|	Gr���%\�j�x��s>s��`H�����<Ʈ�6�X��Kz.�	.S���&��KwҪ��kk��<��u�t�����HLy�����YN��]�d�+qԅ�-�G)Ygۓ����q�X[����G4�Ap1���w��B��O$f�9�-6Z��Q����S���1GV!>�!~w�POĦ�����������+�|mp�f��/�@��)�*�'�����$����Ĉj5�ua�q��/�,�Y�����\l��:�/ PU�j��E|c�bHK������&����㙞��T�D�j�)*��Z��^���gO#�t�7A؛:
�|��F|Ԁ�Ä��C��@)F�n>�ڄ����>����t!��Qw����TԖug�����X����A\�I"�w�tx��D��]V���
�4�1߲��7��h�5kt�o1�@��i��^�����K�\�u9qq�;}eFզ���*�b�6ł�I�i̢(�Cre�`H���pjۜ �@��qe��Q�`i^3�!�V$wS���V���{U�y�� �Zv�<�Y��"h& ض��\��|�{}ɼ3�%���avP���P3H0�Sj�A:�Y�Ȗ�{;ׄ�gO-tO��Nv �ݡ{����_� LϏ-\��XGX�N�"}��t��t�
j�X#�!7�a��o�5J�+���]�۰��:!{}��ۿ��k��vٷZ�-�����>��y��y��w|-�b&.Ī�8�٨�"	�H����b �l$,�G�
>��7ՍF��m���Ȱm�h�_]�_��Pud8h@�~��~T�7�e]�dltHQi��2Z� a�lU�1�<UV9Ȁ�^^�c��wB}/��,�~D�.�$�Za7sR^��uםJ'�cӾ��5`@�:��[�����[�6�x�����|P�& �[W8A=�e�	zz�jX�*~��HJ�
�ozȱQG	�G�X�Q����H��}#�ဖx�ʸ��Z�P�u"
,z\���y�>����mx��\��o6����z4#��ޓ�*a4M�s�xr#���Ø�{yu�"���CL�(��˫��LE�We���ؖ����39�֖�3u�s�YWo��g�j8���P?���׶|�M��c-9���Q��f��e>�?-�#����93�}LNJ���4tT"�����%��x;��M���;lh%t��%b��s���\���=���;2��Î�ﰣ��=�(�	��7���Ǫ�!:���Qs���YY�Es)W�毷���k�
D0��� N�����hk�ʇc��ks�>�� �Xy����`����]�؈�KƗ	����Z����==.�h��`�H M۫h3NK&�O�hOP�X�T�ގ����jM�׍U8_� zA,8Z8˷���}�RA��c���,�s�}�oi���W��-��e|��d�cmפ��]X�i�w
�.�M������e���I�:r�=nx0�w��[���aA"�|_2���v���;Q��O1 MЈYp�?��zA�"T�/�Dbx0��F$**�"V#�D�=LI�I�3N�XC	��@D	yE&�����#�πC��[iy��L;QG��)a��F �v՗�(@�XV�0JI�)�uM ��FB� �E������lЪ����`X�ӗPJ�D[?(o�;:�3L�7���9�O�0
�]C�1���Ֆ=}�	��ӫ��^��R�{��L�t�؂�)�E��k�iH� Y�Ux�
F3$j��u9@Rk2���ޓ��G�%���,)�Ë�S����,���Kie�8��v��Ap�)X���f��d�0��@����N>	�<]?�``��B�ŉᴣ��ܓ{�2K^��m������q��謝B�����L܈�ⶆa�P��߁xo�n^��6��<^���K|���}�݁W?���3�:�TH"8߆h�J�Wy�Tw��[\�?�e��@�w�%]�Tdq��'�QG��i*��ǔ��A�8�QDR���C�n�n�@Cdy�vݸ�%$$�g�\�ʛ�P���<=3�	D<(e���/9���<�(V��}�D2����L��rL���������(��S��2�GX��p2�b�셇�E7�/r��c�Y�f��GI��!L[��o�k�)r��z>�:�/4Y�wuc1��mp(4g�"��W��r.�P��/�M�l�2D��ֿ��EE~�A�+Lc���7��4{��[j����U��84���17�������y���l�l+ڟ`�����
����)"��,���O'��ε�PRo�]��@/W���թ�����?�vq�����sf2�琣�ۄ�v ��@����,�~Y{)���)��C����g6�J�qY�	P�Ы���r����lo�2�ϛ��,Qt�tA{�6����`���彤|@���|��ha���!�AK��h:x��$��$�!q�G����U˙��Մ��2�	�3��f3�K�z`�#;P���dmփ��qڗ�f�����aQ]���c�:���S�k]^�졟��M��P����D�[�B
��b��VY?����a..��-���ׇl�A?�A����0l�A<��2�t�6�}v���3-M�-O�H���.H�ޏ��ʫ��L�'�`B����	�$H�/k�|�k��`�XdJ�VKgL׍
85�����"�Qp����n!zkVV
��j��PО��k/��غ�ۺ�oۺ�2��1&벦������AA�� #<�\�
�b���!� �Q^��yP�f�g�_� �lE6����5�N" �3�o`�E˯"�/§s[?�8�)O��2Dã;ER�Y���R�'��Ƕ��N�R4����Eט8�1�k�3T�'����=���ꀈ���ZZb�kRAX�V���~%���$Mml����`l^lDA��Ht��!���	��͎�0��a�_����+���L=�-m�*��pÙwE�������0>v"����-�U=� ���j�5�ga!�s��)�($�u�z�i��0�����ˡ>=�*}k,��:0��V��d�H?,ʳ�MZ��� ��Y�pUm��:27+V{��w�����.����@/��~�Z�@%�Aѻ KRc�cW�w�ͬh�:�l�Ze(���+x�E�<�&M�8Ɔ���gp�7��y���� �ث���i���3�?׀Wؚ^q�9<y�<M���,�k?���te�7i(�AԲ퀛D){fs�_!��t�+��W���g5��
�=� ocQ!��N�~E�8my:k�Q<>�8������^]�[U��HI��v�ޣ=!c��	k�*-��^���<�:-�KDhg��G�L�|X��R�YB�x��2�#1�L.��E�Oa:�]� B*ߪ���]���h1���U�S� �t�5�`©�:���mEl ��ɫ00{�J�Ʀ��8�)G½k�(y�?����lgr٢�j ��w6;��{�4�L����!iŦ�h��EB@e��x�粷�c�5����5�xY�ph���~�awN�Vy���F���6�H#s�)�!-��(�cւ�O&�eۃ�e�B󭨉�4n#%UUO��`��E�ā�3�u@ �1��p4�U��^S�!ihp���r��;������cҼ���/{v��$]�:�H5��p������Zt�&$힤u�φ�`k�����%��+g��)��v�-R^P�*�����K���;�g�F���<��h�v���[���f�|P�M$�Q����|��@(�0����6�m�>���{�q7��И8Q�Y
.�o���R ��h�Bĵ���st��|�Qb��?��ߘ�{�.hX�=�����(.���::��k�s����[�fE1z���^>�v9=��RQ��/���8g�|��t
���b��@�x�n�����9w�]LY��^�5�iw���*��,���m���q-�RVȖN�W
��3��C�<�/`f\�-C)��qwy�B��Seg��)��q&��Pd���3�S�Em^˚Z��a��8ˌT+z�ĵ�
�h�웠�fod�}�e%�MC��zXմ�����3���֢v#�x^��D�L'�ܼL�-M�n��e{��`he�d���W��'}�����)���V�廤�p-�cy�AZ�*�@�ig���r��y���ǟx�2p���zjq{�/B_�`^�G��!�����AF��a�+�VM����lbx{KRl;���K1+��.�8��6L2��o))ю!���z���Ao>;��\L�X.v�nF=`��"a��X�E���������]xї[ލ8��_sB�K�������Y��̵��U}����D�ƞq0oU���T*�,T��h���,K�z��0�Fw�x��򸾑�qލ2�G�G#��Z�u�r��M�Q�"ybuT[D���x}��5)��I��,vt`�s����'�}��H!�~�&�AƔ���,a`�r��k�1��O��4��.����i�E"]<`������ke�#�X����iZ�����ܠC�\�=j�g��g��.���{�JO�c%��~��%`hԾ7aL���ep�����y7(�
��`'�m�`g��=YF҃Z4(C!�+�g�����/���NC_�d�Y�X<q0��ԵY{����%�h�H�qɿ�K��d7������ś�x>�_p����6�%�qy��=��RQ���Л0�|%�������ƛ�}�/�-;�	E��P}���3ѕ�������u],�>���?GV��_�?�Q���B����n�\�z�%�Z{Z�=��v��^���;���"�W=�&p�\csR'Uy�װy��y[�<7�=tJ#�t���ɍ8��Yq�K�D�(:7�~g��JD��fپ'�,V��|qdG{���[y;Vc��Ʃ��}����U@�76=ӟ�g�#V!�dw�y�����D��kI`le8�u!a����������GZ��R��-��N�՛���"u3<3{�<��QT�Ѭ�.��0
��I^�K%����K+�I��O��� a}��U�1�-�G��E�l1'AW�ʪD8�<�όe�Z��i��,k%��5��=�&���cCќ3���Y�m����ug1�Kw�ԓ\n����#����m�ࡧߔ�A�� fo?	�o�`��>�-ZHru��D��ޫ��J]o�B�T�80|N5�?�	�7��Ej��|�-����&X�a�>�>��ML�@8�,���]�I��ke��K�ȡ�����Au5�4�U1}�Z�z�#;zpB;� ���0�����Kt35�l�����^͚��D�>w�
���3���v͹NсQ	��wF�P#�w)	�?=���o�%x��z����:oYh��6�֛�c
qE5��U�`���2��y��`s��}�E9�~' ]oo�
�֒o��/O����RrʛI|�tXRBҁ���Å	�vhx~L)��[���߾�G:{,�]�.$_�$5xk꜏�q�N���*b�3��I�O�j����R~W��N�E_����@��c�^�ZFϲmS:��5�*�2|.��W�@pL͂q�H�_ݞ�X�"՚����g�1��Yį��F�����ґ⤎X"�;ԗB9Nq��T:��ј�5�r6�J� ��mW�VΝ��V_~���a1� j�
�� Ӟ�G���D��d���<L��'��F^�K	�;s�a�%�  %�vc;�{y
A��a�,�-�K�tZ~bQ�H�"s]yu�Ԫ筂&7��ɻ
ѽ����"�/�f&P:T����]�I-�.��y�P"���t���B\n���#0Y�F3��Ct�϶�AD�{dM���"h&��48�Q�q��s�,b �3OOI_�NK�m�·T����z����mw�2c���	�;�%���s�9�Z $4�+Xg��D94�9�RM4(�Л_��?��3U~�x���J�밅����eb�4�dʀ����;�	�yD����U��(#7��[�(��f؛���
N���9�ԁz�?k��Eބ0U��]H12\�⣔��vf��X���K)�.:͏�7�ka_ӊ#>'G�a�Iǭ`�|n0y;oH��j��"��㎯��v,a���]��N�mc�}� �#W�.���
P���S*��ùD��ũ����rdQx�^�_)s�@��9��:�?�*y9���,�Y'囡��ņL+�ni��k?���O0��9�y�?�^�@q�b&9��4z|ϻ�GW|X����h�^_��7���r�k. �TJ����ke�af�y�̊���ti�,&1���<��Ac�����5��v��o�N�v�WkQ���u�m����*-�ɬUD�˝��`��款C����Q���[.�������rh�Lt�-��w�� 9��dTR�!��%A+�Cڗ]Vْ�B$�fށ��M��)�V+�ua���{��5>N#�Bqee�&��ZH��~Źa�П@��[���
�3�.��xe��;����wwo��)D����8B���{Z��N?:3�h�x3��pn�rC{�TZ
��Fy̍��RD�ϱ�6^�����
hX���P_�,V؝��'���Ʀ�����j$�3;�q���]bȊy]d�\Y��+���n��hq������-�E��c�Bͧd��飼�H�Ƅ&zo�� To��"�g�L,��X�)�Բ
h�gn`H�y��<����GR@։0���+�"î"��P��I
�X��܋�=��0����9%z���y�m���k5Н?�23RG�V`�9,�?�L2/U\����49`f+��ׂ[����tQm��:�J1�9⵪o�S��߲�:���b�AT���ɟ�%w;94�K�"�?EM��q�����4�����6tmx�Mt������2= `�� P�jX^ڈZ* 3k���TDd 5Ԯ��t�S��'v	�ei�|���������VNQ�n@�n���^��=���զ�Ǎ5o��ea�&G��!s���J|����{��)�F�8 (��,�/�?eWhl��ZE8/�v����I�r�}%]o>#((\�*#˪V&{\z��T���%N��Ö���ڱXp� kW|jI�\�0T!���R]���t3`��		C�y�����K�2�A���%7�[��	��ӫ6���;�&Ƴ�& �="(PZ+���\�-���5;nZl�#� ���ٯ2�:��A\9`��5�<�Rjꬻ'�Z+�o�������S>~�K�Pkפ�K���/���q���tހXk� +t�����BSE%�r�[�嵺�S��\��C|�K<�Q��E6�lGT���4N@�SJF.�?�5��<��|j�W#Б��sd�x��r7�)�To	�h��+�'U����ipf�oң:@k.�<��[���F�˙'g��J��{ ��a�\8)/��j�l���-��Kd44�]�	~�e}���gKf��.> >D�t��Wv-;�	�y����B��8����U{#6]����/"}\�f�}��hR��(�̚�w0ye�\�^K�o��-Nk�z�P��F��K'΅��dJ���|@`���V`�&[�
Rw7s��7r��vP��dĺ�Kwa�V��� F:[N���5(��2r��;���fhAa��#�~De�n�?���;
����fU��;@��>I��9�3c"?u��{J�w3rV��+m��)F�i�\�U�@`��MZ�$�l��2X[�-��E�V���⡁/q�ki2 �1�����P_<z\%��<[����
����v��!�h�t�ܐd���S܎`�$Svtkqp�L���e����&�4�1�|ֈ-�v3�db�71;����\ǒHp�zw�3(8�$��Аa���c�B_�w�A�$(���,��׶�hf���})r8�3���f�hu}�~�G7� �7[&^�04�ÆLZP�鄗�[+�Q�G��]?��"�}��u�0L���9�c�{gc�>���3�?�)0�(1u3�� �wsm�7��Z�wb()UA��VNsΈ]��tq�_�g(��j��{x��t�!�WY8�.��G;�����z��|9vo?�p��Fv88ӴFq(��oNNl�*^]��"��޿��nv��"��E��SSm5|"��ĦvT=bv�<���L�i��!1�E����(��]���r�nno�,�Q���g=|�fϧ�؏�U�5�\��0|A׷���YY� ���xVZ�!�@3��;� e�3�ص���Ъc��z�#gi|?O�x��^)�%!6�gO�G�"�n��V�gX��
u�.�v)W�7O�-}�΁ZA?9V����J��rfΩ���B�wqU�?n��F�5jp�it�"y
�fO|�m�R
�Խ�=��������8�Sӕ�0|�er��ዋ��H�u�iJ�X�I���5L-��c�d`�3�2e��^^S�2#�c #n)��"�|�xu��gz{;1�uZ��X��ҭ<_\���)g�D�����@��ո_�)>TA�|��`��L�i+��o�҅����8Xgc�K0��B���컷M�����]��Z��7��Ƙ/�����2$�{B>���ϔ�Бx��/�"���3r��?*�_��Z��e�Eř��� �G����*[�'T������_h�A=�h����������3s
�7�Ӷ�� �\�!4_F��J 	&(6)���K�Ǐ��ْ�Q(F�5᭼�si���g����c����۸�+�'ʗ��^�NpAs�Y�:��Z#E�2m`g3���z��	���P��dMbWCIP�2��Sd�HB���rFnlh�N��]'_��w�טh� ���ݸ�D�B�=�P����\D�E.���`q�2�跴��M�AM�Tp���5�������%�ʪ��C٥#br椊UB� ��a�7/��y9ό�c�zp@Pm�b�/���oT@�ș��55tj[e����%q1V�&�՜���(�����k�rl��}�VٟaAQY>���` �4щʹ��Qr�?���Q\N[¾�(V�� ��,:�o#.�-}bǦ,��,����w-�X��@�t|�E�Y+����]ʬ6�n�w�`={
���R� !��8�'{�����U2\�Bcf��x����������#Q�N �i'�?���ܪT$�	cM��#��h�7f��$8H�B6���\�.������ɒ׽iD���ϯ��Ӊ荃�V��@6d'��v*&��,%��6�9�U%3��*�J5��eȚ�x��[�z�gz;��(��#ܥP�b��C����7��?���q5o(ʹ_����-�V�_X�Q�p�}J������v@�?x����{|���˷wE�S���3S��b�U9�̓Y�P�^Ʀ�&�
�s��n��P�Ow�~1��g2��Z9����,��M�X؞ϚSz�<�Gu%��z��!OMG%r�O*�����;���tߤ����չ���Pu,�����nݡ��r���̈�����2�p(� hP�o��Z�6��r���\bcB���_W�g<��N�3w�ji���{t����Qt��GEv��aVI��1����v�6#�����Y��>�9����ڏP�?��z~{{���������3��������I��@?KL�kǸ3hlrÍe7���ԽM��N��ZY�f��(��l�x�5����.���y%1�G�n�H��J�����
M	��ʛ��&=������
+�+�����.ȓWEjtO��!;jo�i�VO�osC��ʺ�M�\w�?�^6�`Jw�q��J���!z�K>��w6C�XS�HG���ٰ��)�A�XJ�3g�`�������1)w��˒G���ʔ�6��Ė�G�]Q�k"�7,-��o!� p�v��Y�:z�Ae��𩈪��1�/��<��5>Pp�o����!��Υ$A	�L�)j�E[M�1�_\�덌��<�����=eZ�����qB�~^�;O�g���Uwp!J�o��&�k-�#.����r;���ɈtcK��lG�8Xq���5M�YK-���q��̙G�p<A�	��0�{ ��uEZ�/bŗ����*Mͤ22;�w	����k�S K�o�[� M#��� �B�W`f$�z�Q^݅�;95T|��:ŘX��i fZV�n���Ag<���PAiA�]=&��Ɵ�6M�n����Iz��7
RR���O5�ׇ[��$s1����k|����X��_s>FQl�{V9�o$��R�sW#�-Ʋec=��2:�1NT����RD���Ԙ��ٙ\UT1���&P5kX��b+W9��b/�-X9���!}�~}&�
���zMi�8���`����Ф��X\LS��eѸ~���n:�>eT�@� OQZ�
���@0s�?���[�A�괗QS���&~�nD��/��L>[�(��
��1�M|�6FVyA���ݔ��w��X�IO����Ӕ�l�Ϛ}��!����Z	�]�{3,�D �E�c;cn"��&�j���sa���`���?k�q�������@�y�Eg���F����Ќ�Ys��r��efm�h�̭t���<7�6������۔dQ�?:�]VP�W���B�i?������(�>-�p�p=#$�.��ry����j[W�Ī@�C���;>��t��/�(YNz�x���#����Q慄ւ�����\��	�֜��|ǣ�H
B��ɶ���8�O�6b�x�v�f�8���ŧ(3����T�1t��ߠ�fx�Jh�Z���%zc��m6Ӯ�R�C�c�tB��Jz|����������ٝ*7;>��S�īQ^t�Z���oN���,uΗ(ޮ�-�W,��6/<
]����?8��1h�j�L���O׀����,��}@��d�to�5����3=�0���}��i���DUbI�<>b�݇%?��O�"@_����X�;���I/Sݠ�}]y��h�d�x	�ͅ5m;5�����yϱ`�1YV���������|}e�#ۺ��_�D�3�+�mI��zh��˝A�5��Y��o� ��l����7�K�j�������J�.s�5�pQo�DeR��Bc���%����ޟ�����$��U�EM������� w �|'��ʀ�����)Z��N�h�jdi�c��]��χ xZO������:�]��U��J�=5anΐA�ͩ�aB�j���r�s��G)&��D*��2P�C�B��w`�
�Ӯ�2Vk���̆�D}�|��=��Fׯ?��Ա���`8�L���������fs(����33rM2<z)L(S�o���׽���+�w�D�7�<�����CZ�s7Q���)�+%|{��v����mS��,{����O�U��̗���,�z:_H�ꡉty�C��I��OQI)Kh!�:�PU�ʾ hS��֛�n~��%��q���U>D��^����z:�Z ��;}Q�}a1�n��G}튇7D~H�5Xh���x�C�����9��w�v�����.�|�%cr�]�]����>�A>��fD��J�'p�2����O��(�Op���ւ������J-�|SY�zyq��ύ�:�Vx��Y�o����5����6�K����>��{5z'�`p)�L��L����r�u)���R}:��h28��&��'=NJ���ݯ%$��Ba�)�#Ӎ����r!풪%�����K�*������ o+�U�q�0``dw��r�T�lھ�%c��<�]�R9���t��� �G]�R��V�6�+�X�j�nՑ׍����]�њ1�.��͞�p�~oN��y;��>��>�l�GLw�����	'.�ӓF������E|.�kQY�5����d��	�M�ھ�t�c�j��Qi��C�p���J��wO}Ԗ�_j��}��)�_�X͞^MШ����\����./�V�;k{�¾h�g��HDȫ0A��]t��U�2sl"!2䘪�1���
��:N����8|��j.k���'����s�Vw#5?9��u�t|����D'�C�⑺u�h�A(�%�c ;8��1]dTm��hp��e����^���5����9�H�7�wSf�$����@QZZ_���
^v���VO���j�n�7X\r�I�3�݊�sz#���]��P���gc�"���\���n��8�g���?���Eo����J���zv2�:�$��8P�Qyo%������D�Yr��h�-�i�Im�N_��SG��)���'�:���Rhhr�ذ(( �[����	��d��&�7�8���cߩ9�����QH�Q\=��K���d��$pza����s6>����/K���	.���[G �#�c�I�h�%����$��b�3y�+�+�G���Ԃ��$a�r���?^NkeY98ۨ�ŏ�]v�lNLK�d�A��?\�PM�6��ww���Ip'��ݝ�Np����5���K�{���W�Vm�L�>�Ǧ��`�T������(}����b���l�]�N����֜Ϋa&8t�/�I����+ᶾds�����3��[����
��;�;���N���+�̈�R�F��+�jx!�x�o< ĕ�H.Pp� -a��q�>��ۖ`�[�n-ը�,�_�w������;�9sa}�YN���hYٴo�̙9cN����y�/����R 
�ΝT�h����%�m�5T��Ei/��^��<��U�����b������&��~�7�g*X��L�P>��K�I��h��"��z}���_of;<��oC�X�Ar4�9���`jr2�|?��t�P�����|Ůx�mߊhÑ _NF�����\�����z����z'YA2ޥ�u��G1͹�T��R$P���M2u�V��	:}(oc,�R٣�]��a�x�T�B�q�n
9͈@�g�$�ݢu��]��=�����ݚ����T�'WU?���� �ې���.�6���>i�s���4bɚ�z�7��v�U�T" � 3�k(G�Ӿ��&�kn#���Y
��P����h;�w��G�t��� �E�탚)S����?G<���}���e�|�U❗t�	bҎkG�&�U
��<d���`�V<Jb@�%x�k�J�ɼ����A^���;)NH��7ӹl�k��ز.<}
����{� ���Vt�t�ק��󉇟
����_
w7ԾU5ѝvy���H��Ǘ����p腼��N���3� �
�h�X/��tw�4ެڿ��dG4�$k7?��~^t8!�[�L��a�k��"F�����B*0R�,��)Ȑ��Q�u�a��袲PY�R��t�@V 1S��'�(�vZr�L�N��-�o�g�,"�	�e�j��B�ۊ��Sۂ~0@͜�`8�M���>�Ha��E�eTßCg��K�[SA ���'�h�|Z�>8�omwۚL7i&�o��li��mn�z�>L&v(1�ʚ@:�R%�)c����l3��X��rũ���Gk�P���>>�YĦ_��T�@_�F.j9`����^�r@%�Q`��.��ѵ!���+M��\n�c���c&�ˠ^�R�/�$�C�� ��`\�ޣ�{���'��{}�ϐ������\{6�@-���8��|����>�*��������F�5���Ve�h(6ٹ�ĐY�&�@L���8���⨆~�\���.���aC��n�W�B��|26���l�ޞD�����%|>#������ rK�@cGs�x]iN�T6���FA��ɭ��O������E�������dn�ZsjMxV0���]�,Ґ�&����NU_&7a�ݢ��!�&����/�?^.�l�.8}\v���ˠ���ͥ� m��9,�5�Y;�CƦL��|T�#�(�����a��ڈ9<��{�4��eR;�~�);ZT3�ׯb���� �G
�u�3�Ɔ=�u� �r���]�k:�S�y�`�Z2Z�f~�_ێ�h�W���z��,O�Ý��Ew���̳������h�ڿ&�(�eO��gk-*Y!1��ٖ�R*҇F򰴔N
��_'�Y~����K]PR�_�#k�u*K��
yS�?_�f� �2H�x��{9�,"�6��gn����za��Br�)
���M���)�boD�uT�$�T4i�W1DBdt��~if62Ipj�MqB�x	�ټT�\&q�U��4�u�$��..�싮sH���?�AĜ_~I��{�q����V��Y��:r��v3�N�ufÿƒ_?��83Ctns6��=���}��S#�^��,#)fMb6T2��g�euI��Vev1�B�9�Ɵ����%`&ʎ\�Z��-.��,�M�~|���2M%T�1#����3d���g���dc����������Qq�ֹ��pi&!�:�M�r7��1A虌 Ƶ�Ý�����,l�j-���	�P����ǜ��:�Z��͓�<`�"w7�4�_;4n\T��q�yJi�	a(�n�3u�Xn?o��~�M�۝�\!\��jԿWm����}1�Yyk�ܭF�y�E�����Y��r��˟�b�&��(�84�����ZC�ǚ���bӟ�\�`����:���I���M��(_���V/��l2KTT�W�5�@$�(�h�OY���Q�*��J_�C�����MI$`�NDQ�NF�(si�߁Ȱ��,�/�Z���(*2����h��P��°�
��*ۇ�5���C^������@��A����:��q� �!�N��XK�ۅ��	��c�M9 �i!���M=F�mР�a��������Ba�@	��}��p�<��Ŷ���Q
�e�/��� 5ġIa[�cM�\N��
�t �������(?(��Q�/�+��O���0i�'&n�`�bV�]� 6oG�g�oH���l� g���3BE�jq#ږ�����u1�+�1'�p�`���7/��dP:��t�tX?�Qw8�W>�7���K cW���2	�� �Yy�)�q<z�.^�aL�$�G��ԙ�W0R���!@��W�<64���4���(^�Tg�x8�W#���S� d���W"я :M�� �2͹�%��ۄ<tX�x�v�z6�5�� n��$��7�Ǻh57�`h�����v�j�A����q�q3��nY,� ��rc7�jU=A��-:�36y��9�j�Yxy�"q7��0��0��98�����DN���\n�׋��y^T��⁐��)�@�٣�h�����������'�Z�Mqi����P~�N���n��}�9�����@�b�|���rQ��/�fs�qa�ys��L�3F��P�b�[�%{��N�}����z�XY��;��E���{��q���&(��O��MV`FD�޶�{o�2l��xN����x�O�6<�uU��{�����e˟��Ou>'p��}�`9Jiy>=���Z����"!߸����#��D�⿝����m����h1>%�a�ޟ��6�$C;�ھ�� 7P
'8v0m</J�^�W�#'��K�å�X:��o-��Am�5 q1f@�����V���A���Ⅽf� W��'���53V�pX�j[�ǚ�y�H;��(� �!Iwk��4
��ԙ�`bB��}a�����6���]���κ��KM硜�%T��d��u
*k��`ط����Bt�Cy^GlYY�;ᯏ�/oG.O�g�G��N�2��@�'���CG��zn��u͏.ô�]R)�˦�����eca]Q�]�X?��Q��;oJ�.6� Tcr��V�/��t��YU	�Xe��jq��O�ᯞ��yY�0ga����������
�h7QA�Y�-%���!��.7�#�[�\���8�8^P��c۠T�8Ý��d*�T�����ݖ!��\��b�H��}�1^^��U?݆�ubr��`Z_����c��-�m�O�!
�Еￕ*cA�f��QKs'f�[y-�R��> ��Ç	2�U�5�c��~���b��|�)�G�L�����h���-X!�ƒ2n�0{��?$�s���z?'��i�XX]狂��6��e�]�:�.^7�f?lB�p6Z��6(��O�y�)�Ο��f�����p�Ѿ���{��A��Vd�VIvB�%/9i��;鮽t�p�GQ�L���/�)SR5[�������]��Q��S`���S&��뀫����b�5�%�"bMض�Q܁���E���ع��Q���id�!mr�ag}D���X���k��x���?�d�}%�>��"T7�r�A���N���χ�SUG�X~�q�T;�y8xrySD0u��ZG��6}]�=��P�ӳ�+�����;�Dux+	���l_��!
�3������.?W5=+�\�t�6q[��N�9���?�0���v���v?���j��h���j���j�߈�`�W�.stf�/y|�Aq*R�/�'G���9<v��Y��Fi�6�;��&"5;=Н=���_��wژ�	nV�`�'#�O'�VY��߮ZUA�ŌQy|�hu���Z�h�o2����j�N��4�� @��o���&e���'�����}x��b��ꞓ�LPw*^����L�):i���M����;]*�u�$��*3z�7.M�O�ȹS U8Y )2����)O��x�f�E�2+���k��ꔄ^]��ݡE���K�U�&��=� ~J���u���5c���^���ӂJ���6�	����I/<�;+]G�6�Wmq�ko �_s��/��E9���<6NZR'��@ax��ǟEK5Ê�y���dO.������~X�IZď�n��Q����r��;�v�M�{8��͜Ų��1/�K�p����$�痀UY�S��_XL�Ȓ49�zY0����6���F�P$����2��ƛ�QN��Y$/���^l'L�l����^Z�N���	�~
��|#���r!<[ja}|�NV.�ˊ�H��SD���MT�:e�0�O��4&W���]j�^zf>���c�˘������6�( �i�mp#3(��&�O����̈��l)�P����DK�b���
鱃��=��ND�tc>T$��j&{�f4��jB׶�!Kp�����>�Z��v�4sʛ�Zz~ځ:�Y�Q�}��`�|��%�0�9�5���ȷ�d�{Tp�괕j����d�P�.^5]z0#6a�;(xBw�#ͷ&\u"��ڡe�Y��Hg������44�	Z���*I�/�x��%N��傢�w�'����i��	�;�AT^s~�����h�F�Kp��ٸv������GX�%;i�
�ڵ��\ �����]�VP����+��e���l��ͺ�ł�b� �g�
�	m*h����e��sTG&r��-�F�Bĺ%�|5��w��P[�HEJ����ƻzwHU����K�x;�g!�Ì*��ݑ��N���|��h�׬�jB�ྃ���i��3�{q'���o6}��r�,��Q��[jj��*��M�%ԁ�E����� ���C�Ksر5��9Fӻ��He��ޓ��hu�k��bo�͛���|�щ7�.JK�d��N����8����f�H�.�f�B�[/����,Ka(�Bz¯�m5���8ۿY�n�"��&�j]3�k&�b���J�J�W�<Y�%eyI'�3o�$��e�L\�iD1$�}�y����tC>e����k�%:��؇ƴ���_�����ݘ��X>Ƴ��&����r����(��]�^��p����X*�y�.�Ω�q��W�����xE�����W�T"��?��BxT/����d^�x�b�% A	�����`�LA���ب��d��N�DE�\����`��0S�Qf�ƍ�cX��(|���G����U+s��u˾�\F���y7���3WE�]���0�d�gu�M.��J���F�}�J�>��(Y��?=�<��W�����j�ޅ��#�0l~�떜^uPTn��V�
�^��y����]D��o/1���;��Y|���/���I��(q��^��ZGp!/h=��ͬj+�~Z�B�TO�|y�c)Ops��p�%�:�M����%��;��ͫ�L�֔5d�L�������|,|�꩷Fc�!H��/\ډ�7C�̈ǜ��Y���ﱅr��'�ԯ��q�ycl-��?�~2��<���3P��;�whUµYĴ�]E����B�١mM�g+���Wu"�u)l��=Lee�yX9z��##sEY�Lӟ�-���~��54z�c0� z������Ji�����fi������jn��?��$PPz�6t�ĻUO��/����^����׮bMz���ܭ�N���U�fF���i,�.�$�Z��
<�F?�����o��-���}O��퀘嵭�����k�]���6��w��؉��+|^�QCe'M�S�>e2#vі;o��}'c�n�]5�����;1C���^����`�l	T����4mm�؆.mK{
��������I���� �}GHy��r���|9A���N�[
ݳ��8����K��2�e�ڄ�<P�.*�xb�W����Vr���S����]�|k>�r)��Ţ�r�x��.<?̍?��'�x�jƌ��e ����~��I��"�o�H�8.'���۶�����u���c�t�pү�ɐ*��S���;��l�}���lF�+���l�]A��۔�\����۩�_��QVD�������t�Xלs<�/��<�,����Y�~��>xT�����Q��_Oxm/M�����Z����&$����FF�0+�[Nz�7	T�Xv��(X��O�,�3��,=/i����T��xM򺡵XߙTd~-Y~��	��}����uR�
��p�����kl�9�U6�̌x^���-��{>X�Z��Wq4ѸЧ��u�jс���;�E������x��Mh��__
Kz'�,c��wrZ"�`�6�Ƴ7peZ�o�tdeȄ/hkJa�KT~�6�o���7�������ڻ����`�ɿ���J�9������ۅ��۔e1����9-���1���y}�1y-�5����e��e��4���I�C�@��yo�"��G�"��i��O����ҥ\4�ٿָpXN`>�@B/hH3D�.���}r;�5��	��aK��X�Y+ ��*���i1�ݗz�qĮz�8���Tp���n�,��'*�O(T�K\u�
D��%�H4�njuu�֔mU�,r�g۟��Y,��hO�;�B6M_^b�t�g!��;�P��-�z���$�.,>������x*�jzpsD2��T�C���Y:�y��@kUȒ���:��k˹���zd)��ok��t�yW
,.�v���|���ꌐ�����+m[À��*��I����"	�������ލ9�/.;�9R��JӔ�Y㣨�a`+MuyS?|2B�i�9|�K_���XLZe��F����~e�2X)�1mª�b��;����Vg�	]�S8	r�/St��,H��T�e"��-�56W�
��7/��o��[�$�U�(F}\�bL�B���
<B��K!��g���,���-i\� ��!�Jcq�T �w�Ŀ�?�!��\���CCi�Z�,�r�)S�<�����in��P�zw��|�}͈),O6����,�~y0��H������^*���� g
gƑO{2P-����<nЌ�ա������5 Uk���3;GFY$�����7�%!M�h�5�ܗ�5��{LT�*&��Lw�7�&pj�}�ͳ��?�x8�)����-�L����ū���8�j��a�=C�xT+���~� i83J1����)�ҳK� @|��M��I@	�fA��r����S5gHN��z����D��)���0�z
��Q�q*(�D?���~�lV�O��7O�=��K�v[�$����L~�Y�1@D35@}��'��7���? )j����fp��kh��a�Bu��`�<��Iv�����
^>����Kވ򌦗R��1Y�G�T����H�[��Q��~ڵ�d�"�Mh�S�>��cŦ�eE��S7�D��F��+��,�������bie*��?�-�;vw|3�@vO������_�=윲��@��,.=�q�oh���9%I��W�p��w�`�2?��,���^u��.�Bʕ?���n]S�����(�7�G%I��c(�[�Q1�Z��u{{�G�Ν�`[m)(��A̿�&'0��D�����A�+g3O (L����t�V{=����S�d�-,L�h�f���V^�0��V$8�=g�Bt�M�e����?���޳R������>�J�mF����q�Z��n��Q�P6
�<+�{d@ÑF������%�H[�PeW9�'#���]�%�3��c~��&-�S��6�s�A�}9;'�����kr���U����
�0��n71R&��U�TN8����A�ԁ��Y�e<�'��`*�SF��FC.�:e��<��<nd����D����yB��1U�d:�J	�BZ[]>M G��`�z��r�����K�������ҦoW�Ar�m�烱>7p�[��X}����R1��0D~kU
c�C��Y+�����l_M$�Yw4:֙�5��)�Z���A��21c(�`�V�I�5�K^�%�6|��P(S�q�}�-�h6UУ%/G��b6�o���B�z�WA�����&����x�|]�\:��C��Y���ڣ�v�R�B�}k �����:B9Q�C#�v�LnP97K
���ڐ'���	��H� �XL�i�ao��!��}z�,�GK�=��:��3�� �['T��I��
����i�ې���1���PDq'w�@t��1���	����O����Q_�
��%<8��1q͌a�g[�#ƀ�X��ԧ����tE.XCW2��/w2���d_�"E���|�EeNg� �D�ŽD\���]t�!�������]J��Э�j9��u�CK�]��|����
6J��}�m�$-��m�yM%uBT(��6Mtn{܃�XZw�7?���i��)�֎/wBx�p޺�0H-4I��b2�kOI��/�N*\��?���Ew�NB $�`�-Q-�����f��c'j��O�r�+�U�3sj��zT#�5٪�P��Ũ�Å��S��v���*_܎����AN�P3�����l�%ku�]=_;��$�
���z �A�Cn45�� �ǃ�|#*�����J@Ir�O�"��Z�Ѳ���dKC�I某�%�p/|�žJc�L|?u!�� 7�j�	B{Wx>S&g�ɟ��1��#{w�2�c2�-���(�Yy�_X��s����t�jL����0$(�0���5?^4x�M��J��j�})}=cH���kCdK$�-w"�	r�ñv�]j[Bb/�z��Vg̲���8�L�ispk�¦n�L�8)�����h���J ʅ�4��")H�eHX��l��m����L�e������Ӻ�s0��������7�\�B7��
F�C*hރ�����PCg�����]3(����ǉ��8��r2�ڕ�B��bV���6DT�/�=�+�V&NV��@���w��.� �C�Nn��Pִ�b���=L�sZv&����@����C���݉E��d�g?*����"z�K��xg�Î�%��T݅��Ϣ�~ ܎1�/��s�4��ٺ#n��\�G��W.���߱�"��e&'@�Y�Gf'F+�����0������(�gr9�T�Gm�;�{�fG.c�\�N�"j�nn�%!f�������2T3�!0�8��=���Ϛ#tbq58О9c,"5QqbA�S_4'D�M�{!���>�#�8Z�rWn6�<3�]��{��Gf�;|�b���'Fڷ��CB�%���Ɇ�5ﵵ�y��υ�De!n�J#�~��%P�D5��o�� ����g�,f��Qq�Z�t�_��d*���EX8��KhN���K=
\Ծ/s#��#ip^?�������B�G ��(���:xܕ`�:`:v�.��A.��_+S\�a)<�Q��Ԅ��\CG/�}�ق��9�Wf�)"L��� ܲ�X��/��*%TޝZq�߱
@�dq�?ŗm���#��@<�Z��k�kw�g�I(��4>[mݱ����%anY�r}V�V٧���K��@���U�����C��]
D3E��7��T���V���2GBԎ��[86�A�V���..�n�������x�S {-�DG,2��VM�| Mu&����*ȑ��H}�u�n���=&ꐂD�@��ba�K�M"�?a�S���P����0�v�)�w�l)	��a��)�0���u�����K����9�ޮ?|:��U}�x8��}N)���_����D��$��c�|�vzp/��j>��o�[*7R�*�5rT0ᴝ�.�?믔���3V�*����%8VUJ����f���9"�oz�s3m�j���� �{�����������	nI,G���98��fG ,��;�AgMP�=��U��<R'���!�Aȫ�SZv̩�ԔI���1`�l�~h-@s|��R�N�j �C
S�tW ��h�oD��D�=�m�����xz�gơF�"}�G�z��A�|6���R��ۺ�O �wEۘ��_�����i�n PL�&���R�^�=��?�*j~@"	0�UV�WB�6ħ}+����)�b_8�6�� \r���>��v����,y��%'n�W��z(kh@(��ť]�{�'��g��I��j<A		}����`�u�S��Mn3����s��&�E05MӰS#�F#�YLxdi�i�s�#�w�|z�0�&7�NPA�5Žߤ�����qy��k��}������2UtV�J���֣V�d�U6������˔������.���2�Ƕ#7�c��EO!ӛnlkty��k@`]�q�d2fF��(}����ʡWxu��O���EjyӃ�|
���R�P�%o'�Eܝ���}��{v��1a���}��P���(�W�Կ�۪�Ѝ�ܖsmM�q����$��V}�Z����c���Ыv��P���\(q�L�W��U;/Kq}�����vb��#���3ި�Y$A����+�U�򜣆�����P��7j+���Z`*?G]�;�V�!%�{p�ޭc�]AA1*�ڍ�op�՛��+����!7xD�<�w1޵�p��K��z�����.0
=�7&{H��n��IS��s���=/g۽r��8���������.vC�и#�	���+[�=��jqC��(�#3:�aB�B�����Vj&����6��^&QM�T�ϥ"b����Yg1T5T�Ŕ8XO�EP��m��b��r�)O	6��X!����A\Y�6�f�(��k�Y�a�oY��"�M�X~�Z!���}�w�	n�V'��� �r\��Z7����vzƴ)!��6��aN�L�N��zI~�����z��ٯ�ub���fDaBX��;C�@���-�f�^sbw�ۇS[,�ޚ!-%��5O$����,j�y��#Pn����#��0�K�$�Go]n�]gi�}o �*4�ܟ�I���S���c�88�]�4���L��	��?�|)B�q��*5Ǝ���b �JUR`���]]�7��[_Β��!�)��4��������w�s���*8���m�b9����������K��W��kl�ڞ��=�ia�X����tfkjB������u�����y2L��cߣ�uZ��'i�e҃�r���f�~K��a}��5(��H�����w�3���!�H#2?L�&T��rw�p�Q��LBB8PKݤ�L#��
�Bf}�Y���˷��A|1�4�mw��w�:ѷD�g��͑�.7�������Kn/Ab���a��)5J\P%8e��c�d닯@�.�2 �]���8g4n=N(J��\�]s$\|I�<��B����\J���"G0�ln։v18���s&�^��������ڄ� Ot9w"9n��苽���c�Oޚ���Cu� c�v�B8&B�0!ב9��~��^��_�q�Z9�ü�6HY�2Z�Z8��:,'м�q4�d������)z�"���W^��C��(������o_[��E3�uiב�k���A>B���v�R����i��Җ�װ}�6~���u�����:�OG8cwtQ��\�T={ʬ���>���D?����3Ӳ�:A/+�q���֭j�\���a�t�n�z
�L��Fi��O����kԃ����������AL�E������nO�ܑ=��ҕ���u݆`����,��yǝh�G���:P$H�T�,��hr	��>P1�j���тe(���F�x)��x-�N�{��~R� @K$�sR0�MJ�8�ǆ�@7e��c�"��LØ� �.�k����@��Y9�&%@����w����:��S������]Xkt�Xl��:"�<�<�z���}�vdd:��nl�Om��2�v�E����<����eGh�u)Ռ�����n����R�w-�w�%��RJ�䲥\�|���x�W_u���o�;W�4��� ˃� (���	��ghG��@�]P�����z�2�8=��xyW�?�R<95�[�+ڋ����_��s���q�}z4q� X	��5TP���������	�q���F��1����K�+	A�q������͛�0S��1C@���5^9�T#��ۇ$���!���3���s���8tn:�v�k����˴r"��ͧ���ϊy%;��,���ozB��D1n:K�L���N����b�q����-Y�EP�#��1w�=O��Of�u+)���n����ǎ8�=����_S��r����,�Ӳ.��:Oڝ�m���F�I,c�@�|�$4%I�����`U1���׻t��|�ھ+�̥=�@&<2��v�/:���| ����^�3����; ]ͪ��<�b����3���^�����xL�`d�r��c:�9Wg9ƥ��FQ��M�	NB��~+�����ig�;�-Sj&��^�x�}n2(���=;�(�v�%^o��X�$����S��=��7��@.ݜ��RL���m�jG+z ��i�Х�$\�B7����s�@���5�׌��|3��G����,���>R�^����ł�A�*gh;�S�iP>�KCy\3��q�Y �2��T�@��}�a_�!ۛ�t/��<�ܝ�:滄s
iLn5��-5��FP�v#�HN�I� �����Vxw��i�`��²<�'�+��m�EÚB�<9b�ऑ�c����`yW��"/���$�β�Z<v��.�mVX��A%!REk�n@2�Ab"A�#�<��2^�^[��d ���O������ڸQĶ�UΛ��	���p�ݼv��������0����B+���F9Ll�8L�6����#32��oU_A�
�w�1�m�04$��;�篞v�GP �'V|3rp�����^�*��16�_�!����5�%�t���+~",���pQ�g3�ytE�E�"'�\�Ѹ#�A��qю6dJ��K؜Y�-LTgꧣ��)j�Q�/㱣f��}�
�_�o�z��ۘG
�u�dĹ�β���bێ��wo�Ce+�O#�������>�͍�Y+Z@�nB��$yL�-�FM��|��D>@�F�O���bW�ڔ�g��)�.[�ZF�.��7nù
��|%�p��9�vz�>���V7ӵ$��t�������ɀ���ψ���2y7MY�!�((����'�曅 �����t�����y���eE� 9����*>�R�M.�-�B#Kа��i��d�y*�Đj�b$���
���|3aF��G�l8��@�{j��z&X*� ��[9��P��
��~/�/��<�� HL���W�9X����<P�P�������.q��G@�I�jr\���|���n��j��?��1�V'}�C
�C@�1=��06��
����W�v*e�;҂з��-pr�i�;�o5��ey}���-�>@T�k�p����
����V?�ّ����124A��ڣ7y�ە	��c` T	3&��!��G�#��p<���P�������M}Iq $���f�*�6C$-����O��`�OܜI�vyk��tc��+��ܸ�X�v�����+�ҒR}A���1,�8'����T��?(�~Z_K�j�����X	p;
k �>�ǕږlL��0�j;���Q[8����G�2������ S��NAVR�<�����
����y�7n�5c��+W4<��b�ٌ�=mK� ��0�ҴЂ��BR���_�T��>б�a�X��Qg�괔���Db�K�@<3l���6T����YQ�2	��g��ĥ��K
���v:�g:~����j�l5�>C5�ﳬ�����oij��Rl�l�i�p�y��L����^���}�L���d�Ӏ<7~��b�<Y���t�xT
��uC-�Y:y�QT�<�X�`��7/�L��d�?�GXL�|f	p���P��m���z�7�VfҸ�b�=���c���`_��xr��H�po�+l���i���ޚ���XH=�C�_t��D�cP����.�BMM�J�����aO���,3�+
��7YW�F0L4gn��;��
c
n-0*��xTC3	f���I�x �=m��\�|�� l&J���/v������֗������>�a��/���2��A���jВ��
~ �F�8��h~�C>8mu�a���t�Y~Q�q8nPq��A���	�G���A�hŊ91��;�����~(���:F[���^ۯ�A(*~��CЁ`3��3-����u�Et��kA���I:�C�wE@��m�vaiv��:gv<	�vFu���8k;�ݹF�u��c���GV�iJ��v��a�e��?��aM���0��ޛ���iV����
�zh�U���SUQ�5���b8�P���Ga�l��@菕��=�a�T]=��r���3awww��f�g���;�Ƣ����:������b�>3����g,n�hʆ<nԇ;ԉ�;����q���/	2�̰P9^���5�Y��A<� ���wA�,���6����/�74>O39�5��0$^|ߨ�y)>o���E���f�'��ۨ�bZ�h��C���{r��P�� ���b�yl��{�^�� >��7�ׅ�����f��qes�G%p��mGp �6v�TYY��M�������dw��|J�!')��|�zP[�����d��/)y�诣���DE�_F��R6~:����`���CU�m�Ŀx��.O�'��B���>J�]�]<�ĖO��J�	��f�kJ�E;�i�� 	�W��B/��D_�x�.Z�km7��۵��rVI���\U`�(�O���|�[��/6EV=�+��v��%���ܢ8`L�+�#BR�1zZ �"T�I~q��8!�5V��pi��38q��T�Z��Dr)���Q���s���܃�+m^\yt-×�lT�ч�3�|ot8ZR5�bn	2�%`��04�d�aB^4��{���U�T�Y�,�E�S�P?�/G�&��iq���j��	C$H�!*��s?P2Wr2vr�n3��C��SX���A�ik��F0�R�� ���)����G�Oh͑b�&��k��ς��E���Hg��H8
O��Y��a@��� ��j���C` �B��TJ�%��I���$�q�Oh�K
���?!��Nh�?�B�����{��܅d��Z��-
+#q �y�s�Phm���a)�`?��y�?��OB�lSޏ���s�&*}�5t�w��"��?�AS$�!���|�i������[D�jw����?6���UW�̟���k�L�`�����CR�[42h�h���Cⶅ?�R��2�5$��!3����ꚊH��G��(&�&��j�'f�)#K�-�&!���B��p�8P�~l�����~� u�"r��\�ȝ���z�B��7��JU	���5'�v�[ag��ߠ����
Q� �A�4�R�!'i�Qg�p�� Ɏԇz�N`i��Y�d�Kի�Iq'�P���M��Wq5�EC�P ����H�
�C/Ifx9�ǒ,V?@���=�?J-�\�>ް"�b�'� ���5�(���c=)zڪߢs�A�̜t�(XQ�4H�Ұ�����2��-� �=DtRf60K������#�}H
�M]i�/��|���߫�������n]iW�}�	_��t���,l��b�= c�+/L��0�!,K�� �� �H*��hPj����J_���s����M:�&ް�[0��A�x ů��6V�ǩ�7���Ö;�o/ w��/2��#�#��)����%W:��$5I1��(j�!���Q�@��$�u=��?���j����u����\l �o���l�+�
������T1�� ���ΰ���Z��[���_]�v���o�3��z���(*�@�L]%a7vR��*�;���7K;��}�ӹ��~)�R�c��[�W�WB�4[f�'��*QE�q�[�(wȮ���#�ז=�������v�7��TV�����:@�����(df��ޔ��Y{���๸~��p�z�y��+�avG�4�U���!��-����j�]��dg�>�B�Sbu�=>ڠ�>\��j1PY}���2u��;#u�쑞��<�:�x���q�:���l�Wj%R�{x[�^�ȃ�A�n�Dl�|��<��%O��\��u���6I���8$!��L�J�щ����u�_����o�}#<}}& )G�òT�H�q����ڞ��|2R�]�3�!��|����g����(Dc���!�	��q�ߗ�h���N�t�/�'�����EB�� �I�����&�T�5�(f���P��"�B4Ht��P�:25��ȅj�#�M�~�^��ܱ(��NC*��N-S5�&����;�m�������f��[w.�~~p�(�����ŏ�����3��A�;l�x�{Ux�zg�\ʱ�%�g ���}�O6��B���M_�?Q�������[t0
����PT4a�hڔ���������oF�2rrv�ԛ�㯅^�q���Ǔ�����j��ڼ	��t�HE�ނҫ�J��(@jD�H(]@�H��.U�-�*z��]��7�f��53��䞳���쳟��uW��E<��J%�И����rC%6dA��{�f��1�E�5m���_ד��Y�7�����)��B]g�O�b/��)���yy�&�4bƋ~U�Hs��uE��inl(���L�jt��`��N��ht��n�P����W���a�雥w�~�JV:���m;%�mB"���R ��{=߾�,���r����7����c�V�,kC�rw(*�e���#���v�F֜�
���^	��g�?:bu��;&Ism�U�f�Tf�fZ|�]ay X�3����>���޹���Ns<�H�d�@�m�s��Ϻ>���|�~���i�5%�s�hc�k?T�v���eH�N\�0ְ�[�im������6L�!�$,Z��ɋ�f�V06}��S	��3�,�q',���:��jģ��#���J��?j>3��_B��t��*�h1{�yI	���T�ߏ��2�kJ�"�\O������_�81r�k>=X}�C�)��>J\g�	H-2L��#�`�V�IǟCIqd����!��6����x�X1�8�*���1�dE� ���^���X�J�"��p-�N^��*��%l�_��ʇeo�^�to2<�����uRVs����\�[qO���m�̗��>>2ҿ���P�g>�&�(�_���d�/�Y��0ik	g���)�
<<c���A᎟-��L�����_{��tv�����;�/R%{��^��ף>�U��W�,���"�3d�{�²�?,9�5�Ɏ��
�O��̴�&j�[/�J~���ݏd�-2"�ʌL��#���X\��~�M�W�-r�#࣏Qq���VT"զ���d���h�R9@R���ё��ExDu�u�?�ѠN��9f-''��>�6��Bt z��ӫ�(�
��틮Y�AKE���.���鞲֡��@k�U?V�Zd1�2�$wW�-d�@&�A�\���A���hSI'T��C�x����&�NN������IE4V��J��JD�Pxj�7�8�^[�t���%:��!Q;NO����;��@��X�FQ {�-�w]p8ִ"�f��[mS�jW�l��Y��#��4O�����j��
��g^T�s�Ʋr�u0��7�\�Օs?|��u��������f5�Qt�E���OP^O+TY�k{~4�|
�#㝬��M����p~��HT�e�_��V4����'��g\N���J�|��do���*pNnnL'038GR㆖�s��o������������+/(Rh��z��Z67_21���6��5X�̙�݁�#�y�@D���P1���@���� ���%��a�D	Gwd�EX�)�1�/SMw;�>��Ԋ���=LS��[��P+ d�95� ����Ŭ��z�k�U9'�0KY�hW �Z).Z_��?�h-�D
�BRr��L���q���n:G˦*"���
XSu���%�����nB����o������_�#Da>�A����(h��e��J\,��E��"�ח�>0+��o �#�[�q��B9�Z������ 0䥮W�*�!����;Z��@�:�O�@P�m��y�0� l�#�/�0U�DH�Y�E�_t.#?T{Z�V�L֗��9�1*��;i�0�m�����'�̽�<v�T�ޢ���/4Є�Z���J��Vkf9����FI�T�ԙ]Q�0B��N���{!�6q�vƻ�
��O��C�R8�����Z�	�Hۗ�u|����"BZ頚r��i�v����ɩ�&���`��:c���mK�0 �},��ϖ�8m�|����a�ʳ�'q��$�W�RG2��&���;�|}��� ����r6��J �X�2$�����R<���!V�a��PI���{M�Fu�٫�04��+�\��7� �_Ri����*u����'�Y�,���"�Yp��p~��6vvvi))���S6�2>Lm�w�2���)����2�2R����<S'H�T�d�
lsC5�4��?<�6���`?+�4�(X_�[�l�k�iZq�Jz�V;!z&�+�����m-�2Rl=a����𺵦'S��9R��btuQ�t��9�/u|"lgR'�Z���_�±�+V�8�D�h%\W��乚&�7�mJ$���;#y��O�z^x_ 8��y{���ADa������.��x=���D_��*+T���07�5e:��>N��(�][�˾8��ୗ;D��0�����Y�8����[�˞9�����q��G���b�ǡ��2t6�<т��`����x���v�>R)�k����'���/����#d={��m�Y	~�b#t�h,��.NK�V�+y�YC��.w�NYT�kI��>��E�)�-�gJ�.Q��B:BHG7��n�s�����/^�s�].��;�@�Ҳ��g����Lwr�H}	�1�� 9fC
}@5�}��i^C�^�V���q�#�9�U��a��~�O?�
jw���\��&%��z�	�`�$' u��:�k.^�׹��{��>�_wڦ#*���_��g-Q~Q�2��E������z�m������"�$�S�|�E?�h\���1�z*���.�c]?\]s:k�J�/,P���S3�_�����_�ƪrEB��K��}&sR� )i�Fx-q��N=D����!AEت�il5�Fh�=�[͜/`�k®�xX
���7�0c>-�{��L���[��m;s�S���RHŠYg{�۷��0�������t?�6�n ���X5U����&���n<��u�r�JH3ou�˭wM��r��%<=+7�C�ۮ�Q����rj��T�|��Y)�N���*z���Wz��Ol�}�~6��W�L�2�{����j���(�d�HY0N� ����C�ng"�Ķ��iХ����j*��ZFfl�	�C_��n��A�6�"$5��!�K�1�z��)�;z%�^qj����b�w=��d�W9]��<N��.�,Y�?N�n.������O�"��3�fl�B����.�2*$���T�g̕/�v_J��?�jI,[e��{w-kǿ�p`���t��H�ÖN�p�m�g9܂-F��2��8�b�M��� �ꛗb���չW�'5ԛ�NW�P�̖y��&j����p�7��p85���[r��$8�֔~0NC���H��k쫇a|�yee�1����'F�]+"�x#��zJir��b�u�CS@06��4u�*Y+�	.��'��ƦE�VO����^]�*C�{2#cS<X�Ɔ�j����w&s���Vz��eE�R6X��F5�g�BU�t)۔}��0{�)�&p�,WEP�tɧ���MV$�΍�2u�8�������\��;�1��𫡌f�J� =�ɒ��w3���W;�M�b�*)��H��W~�V�I�5�O�{���;qx��o��P��锃"����	�A���Ch��*�w�Zݭ�^�O\��dx�i5�;ٛo�ہ�q_����Ę�N{�;���h�W.V0�x��"�v*��ʹO�5n�������Y��	/Y,��7���ke��A��ƎW�]�7��/��)f�Z�X	��ɭ��5�"�j����Ki��fY2D5�ۯTm<v��&=ӝA�m����cU���y#�c��8�O{�^w $��l{�@Hh��0�o�k>و~����2gH+[YY=m!��}n��m�7��F[6�D
�Gp�k�/�Z����ܳ��YJr���8U����rwj�b=cyw�i�����qc�˾��?Dpu2��JC��M.��ޭcA惱�ic0_����+�_���b\g6��:_SC.�,���!Q�]''��i�#��n����>i%���L�%-A4�����V^'L��<"\��saw탹��_��>/,^Y`�:��069���Zu�5;[AA��<X�#:��<s�������#c�����W^R���~uV%�O!
�j��K]$�>i�d�U?z^�����Y=�[N�RP�?ٞ���޾�>:�w�Jq�i��	�\b�����������[bbLKU`1`�v��[��z�ּ��\���N3�f�������sۛ����k��V�_(���N�a/i�~mZ��^h�x ���;�7�[��(�4���s�����M�;�g>n���舎�6��(�0���Q,>�/l�HP��!��3ȁ��� 1��}�Oӕ������L�Sp�w��چΩ��HK��r~�_��{tyZ�`�5f���Kw,�(��<C-�ߺ��.:�Ye̲C����D��$Q]^Y1��(�r���Jng��m�"�5�������ۘ�W0�Ǆ��{���_cA��G��xm��g��M{�n��o�6m��ķǊ�o�$�:e~�.6m�k�8f��g�����T��"�U�&�I7,��t��M�n��C�񍤢߷��'���ȘE(���}���jK3L�rk���A��D@���ag�<eD::J�9.]z���%W�֒�O�H�̘�1餛a;�^����5*�W�I'����JR#9�@W86��tz1�B��!��H�9:.�R�`�+���n���L��r8>"G�!��Ǐ2����F�`]�]gQ�4����ɻk�$��o۟X����{�L���./��~���ߙl
�%�������?8`D
l�I։���Yg�8�����RF��U�8�ň���{M�z�6y�vZ��b�X��;e:)I���?=��o���eⳁ��3(�Ţ�$��{��K,W��fw�d���v��@���g�B�s�㙂�tl<QT@;�~7gw�������V����;�� ���lHK���,�TΘ��f, m������,�=f��y����	�I�m����ӂ��Cb��	\?��E����_��ֿ��.{��������Pq/5.�����Z-G?EQ�	1�%�@ �0�):~�w��d�h��#f��Y��4���<fox�D������b�V�"E������&o�E���jT�b\Z������r�]32���E��-�BCp�������&�E<Id}���"Ƴ���6lT��K�z�ļ���;�4�7n\|��[�J�lp���!�AD�x��0Τ/K��歭�­:�8�+]���ɼ���J�Q 2��]��~��
�)���x�`��D�00��8���/p��^��q�ڲNu��[��{-�2��E�j��y��U�J$<+ #�VW=�q�&�Z��Y �6[�{U.Hd����%kve1���.�,z^������%�'���O��7c���H�+��·}��㶞
��ށ˖hj�ӄ#��.o֯tZR|�k�/��)#y�f��'�H@fXs��n�Ш"V��m��*�U�ٌ�~�p',����~:�\?��P���������\+p�gkP���
@�Z	��;��Ջ���@(����d::���)�R/�v��F�6m'\ھGt�q\���3�;��~�0�Dt�ot��t�ԁ���ͯ��q�r�p�M�H�g��d�~���Jf�/#/���a��ebhg;.�N��r��͠���p��޻�$.ζ��NR0\;�hbi�>��T['B���Є"�6!M�SS`��~�(����z(̋�)�Q����D,7G����`���o��JUN�GƦ��`;S�/XOqY|=gr-ѻ�N��!!*qz5�^k��9ĩ[#3(Ʉ[�8�����?b��K�<Q�$Ԟ:B�n��2�Mv�y����c%R�nL�y
�5Z��w�/菑��!/�7*y0���*�:�]������rtŚh$��ܸ�I`N
�K�n֍�t{ᒧ�e2�����K6NrzM;@�-*��ǭb`y�^�G_��[�_�7jj��1B��c���N0�V	���b/A%^9���y	�r�}`�t�w!�C&�|L�y����ߕ*Я:j�O�@0rF������(��R$�dg���x��S�A>���ڄ��y��������:Ij�ih���c���:hJ��Dm��G\���3�=�F��?b�����������Q��d7:XxCj���9N������(�H�-�%���?x�S��^���< eK��q3�%�e�(+��P>=zs�E�7Y������,�P��P�Y�*��2J�~��DaT�=Yb�m�ű��������� �(6Q«�י?�싴yް�[�˒Q��<ojoh���P���o,����!x��E��k�o1s�n���m�&ry��;s�KZ��"P׶���2UK�7,��.�~�&˫�I qs�QOV�����)�F������;���51���[�G�������6��Џ?��i�W�~/��%������~�,�6pus���fY�	:"�jl�7���7ǈͻ��G�������.���ً���<����`ff@�����!�G[!��� �t�lοi�إ��C�8e�6��g+G "�� N��W��d ��i 0 `M���i�E����n�mԄ .g���w�e�� � ��u����3 �\�Nˑ!�/{ĭ3S@3/�T�T�~������`�E0fi�ׁ�~�гF�6ZV ����|h��xuۙ��; x?S�n�O+d�%hX(�U �
=��]�A���b�
���W���+��
`y��%7�؉������"H��\���V_pOCf���JNoK�!��ED�Q��2�j��z��w�h�|��O�ue�և·�=?[�UC�R�r�=�a��+�.'

�Oߧ�A�>�������+&�����D�C�+1�\֩%�������ww�G���G>���_og���������;��D�큸����������޳����U�n?�/PK   SH�X?S��� 2� /   images/99226213-8268-43da-ade8-d9d07cfcec9f.png�gP�Y�6�3�3
(���J�80�d$g��AR��!I�,y�$9i����LJ݄&������y���s��rW98���k�u�k]k�C���.�\B d2O�VA H���$��̓�_~u��Q#�7��+��w|��@�� ���f��
|󆋔�������DrX��8�<w4�pp�Hŉ� �2��架������ge8p����9~�����9~�����9~�����9����D�a �6a����s�?���s�?���s�?���s��W��
?���|���t�+�p�����q��ds���,�r3�A���7��vaj�(��%'�	�ψk���XRKj�^ی�����~��Gz�޼nq�"�s�lz�c��*'��B���G��*����'�t�����Ð����9~�����9~���Fy\G!�~���AN{�8�֤�M�,�-�U���0/��w�Dd�-�h/j�`��z���L��qe%eP�Td6�`�$!{+m��+�H�0/0�EV\&.1����2wV�6Rer��t��=	���n8X|��^�V����ϕ���-¯%> 6#�
{q�$-��6ﺴGDW`�3�O�5wr�~�;�VNYv���.�7N''kg���}��:�w4&vy
|�4;�k��:�[�$���L�Su��u�w�4���Yz�+�,$d1<�nە��f�=*�����o-;+�s߾k9�����#����0I3��\�#n�-�1�i2E�=�]KeS�g�~Q���z?K\���N}��N.'�M��x)~M�銶w�����2�-#�z!C�܁�����k�U�<K���5,Oz-�e"l�k�xͦ�ٻ��Ǐ�U2�+u�D��uLǭ?U����{3Go}�5$H��67�Ck�g0܆�����<�s���?H�&�����i��rJ=��k���p��ҁ�Ɇ߿Q!aYP+ڭ�ұc�����X�."ί�b��$��f�@�ى�a>�[O��w ��[� _7+�����~g�EG�+�}X��$�qf��q�VB�<��C�����B�o����Y�xj������g�bh����>�ޓ�̧NLPK���ߨq�nd�����B�[F,���O����o��)<�j3����J�-�}^3�S����q�o�'<}'�0M�F��`7�bqmwi���~3��քQ���dFK[XQ�����5����b&��-wd����^H8c�V�g=m$�,�l~��"\D������ӕ-��/Cny6�*�)�O�|�����8�??~ZK��ɳ����[rm�2�#i_j>���1wY��l�[8W.5���P��D#熆�L<������"����Q]��]s��蕄\�y"���;�˰��G�v$��T��Zۭ*H_ݥ��<�>�e�g���P~8FoY"4���i�ɚ
�29�
��g�'٘,�����%|�}��ݙ�F�k&�{ټ
/���\�.���� B�v�ώwt�m.���v���2Ln�E;�3&�e��Y�zDU0�GѷX��R�޺f�&�]0x�;S��>	,	M;R�v�-�)�Z?3����Q��Hs��H����
�y�٩3摝je��4���%{c��E�[::4j���T�/��~)0���o lC�{�݌$O�4{!0uUe���1c6�s��a]�Z�~{0�X�����,��M�4-�F���z����;�N<"O�?�4�q��|�ɗ��Z�+у���[��*�������^�Q7�~����w�㔭�S'����:�X�,�����������K�b/~0
آ����nXn��z><Sj*<�Ij���}{��J��⃖��.���C�\�r�J�l��2�|�-5��u�I�>6k:��y`޸?-3��׺8;K�{�H��d���A���G˝�����ȩ>�ZhO4�h!5n]b�ݫ���R�4�W<+�Ej��7i��BS9n��;xZ%�	?�8 s�<n�%̝oz���(��-��J��/��jX7Z�����(i �_N��Z�û����y�soձ1w�7������2UOZH�N�-�Z�G�(6���oEuE'�pu0�*�S?�=_B����"�/FW=����ټ�*x'D}�}�6�
�����u�:�j��:�lГH7���3Hk��?V{�X�pEn9p�-g1���a �������5��!S'�[ԗ��<`uy��mZ����ݣ�<n�LKǳb��c��`Y�4=�t��?�����>n�~=�-?�1	�/s`|��R���x�g��i[k�����h����__�J�U:ڀ�z�L܃��._{�(�%'^�� �N�c�e�ڔ>���©��3p�B;�,����L�:6h�z���"�Qy�*��hu7r+�Z���y�6��s���Rv����Մ��eܹn���Y�ۏ&�>��[M�L�T	8��J��q>�x�%�ɦ�lx;��ƙY� �ZR�pf�u=wR>�:	��l\�����������(����`!�x����s�Z5� _*�ȩ��@�a�=v�0]��0�-�7�;��ձ�i�&�6_���<�Ik+����>fͨ��ѵ�N0CBK��R��J���j�u�X�N����{���R�6��t����`�g	nK�3rT]ݝ��B��6�|1��`Ba����9Ob9o4Bz�5b�V>3�s� �8	�c{7?�� ύ�b��.�l�*_����N�6�~?y���nTy�/~�8,'i<#��Q�n)��������h��ܖ���7��}��c�:z{��$6N�����:���g7ŎU4���4�}	M�M��f�5�����S��+��pz�e�� 9��BEؑ��#�*@hL�N��o���M'���E�e��h��$����0!���d����}) n�+�~�D�is�=`x�� ���q��$ bƱb��4���/9�0��������`6�������e-w��俀��� Ä1Koc�r�o�v�T"5>������?v� @(zP,{��9�/Yw9f�k�:ͭ�V��H�}��9�Y�o9Z�t��=� ��q ���[}�0
)���|���� X�E�������ѵ������M���Av, +J�X�<>��zFk`jF!(o�ӻ�U_;�����6}�`�p�=�5��e��������؊w���ǡ�����&����'W�Yɚ�HI�:r�������������Իk�oR�k�[	lJXN(a݃���-�������_<V��(��Ow�f�b��g~���ٗ�޷o�h��j�����铆�R�+k���)E��0�GwU׫��<�ݹ���Yh���.Gu>gx��l/���u��j�$y��h�����S�gE D������i@�V,�(��8,=be)���]i_Q�˸��|�FO�������1��U\�>ơ6t,��<;]�i���C�&?z~>%f����V�_���x�f+�,�`�����A`%���Iك~�llZ(/4��\g*�}�~�a]#�1�IK�
�o�z��bAz����P���}ε��1IŠEUUt��1:���0�{Ӿb�=�N��@��[������^4�7r�?H8qpߺ�yZ������s����~�y.�~�y�h� ���!~�2���0�����a&P�so�!l�;qp5	�RPW�hN�>���Bad4ڴ�h4�%ho��r�Ǔ~�}��ܼA������~NGǉi�_x��	C�����  �n"���P��;�Y�th�ԉ����M�!s��y[�y� ��2ǬK���CKF�4�f���ɾ
/��Ryp�`���t���!3��z�{F�Q\�[o�h�(�A��&@�h�*��E����U\��Hvѫ��Qx��0W���z��7!��$t��2���,�mO�����xj�ǋ���p��q=��_��7j�
���S� b��o����@�[�_j��(o8Z�W1 ?"�4#��ɉ	�)�Y��E��<��f>͝�M(-���}����E]u����&�j>��b�}�h�`�r��*� ���~�
dG[���s����'{k�����hvPO��L��_����/z��O�	��wK�D0�P\R����=S*���Mx�vh1C�cܑ��U������z �
 ���Wx����ܽ��aGn�s
��P� �����@���Z1��{x���+.~0>�[ ���큖Ԝ�jWGwynˏYC���ì+��֎������<����jEmX^�J�����d!�kEE-��������A~QD8F���İw�&~�p.��B�� jͬx��� q��E2�@S���Z� q�1sv�t���+,m�@���l~�5{�R|��� U@|��40?��m������F�O��f���:���pi��+0G����$`�ׂ��g���Ϋ���>R�Y�U_���om�MT�xy���]��;=;+�� %Y0fqiCܱ�>A����V�<��P��3�7�mf��w����pg��j�@�i���a��R|�R�0����hh�2�����_w��f����������Oq
A�j�a{l��������}PB�~`w�>��&��(��R}þ�E����o�9�X m%�s+�F�����ڽ���%q`�y���S����9�$����i/F0U��g{���O=�٣�;�^a��SBR�pt�cݛ �d���[����ef9�KA�v
��\��|�̜$�JN��N~u|�k���\�6�d�/�1fTpxog�2���?���'0]��z_[hId�߯:K!\����%8����}|/��FV ��((�~��rV�ӓʏ�x1�A�ܪq�ַ��Ԕy����� J��R�eT��m�~�ǡl����D8��\ЃY���}����;9��}�rR�ܷRR	3ƒmͧ{��8� �(��*��XD��b��2K��z�
���ݵuK˃�)�Qî~ȩ�PNh���M�,)e4��+����gp�X.xtd"��U�gS�xmخ���%Ey����ۇ����ع�����)c@��r�?{�TlH���Fn�U8CFf���������!w��|#���(p�7�x�b��6�ii��}6����b��?tG��g�K�R3+�or� ?d�G^��2�e'}5��Yb���s��+�_������5��ܤDV9�P�ׯ����^�

��3��ׄ!Tφ@A{5�E]S_EP��GH�l��%��a�y� ��#���L��RT�-�X2$ز�L�ҧg��Z9m���D�\�J�+�rO�ijJ����I>-��y֕R��1�#��s��j�"�饻�FoP��9�*e�F��{}O&vd�ؖ���] ���<a�%'���FFJ|#(��\���-���XcU
�{m�.|�Fn��@���:`;��߂!�:�$��I��-����{�	�+BQ*%O{��N��d}��K	�����(��r�������}��`���6B'��rV�FYv�w-u��adх����ވ}F:&9"R?��@];�X���rb�SW��>��'h���Us��M6��i!Q��oS{9ʖ������?,rUPȴ_YK��Q�QZ�����ҽ��d�cc	2��]�ZZ*		�q��^�k#>�xlE'�
��TyN�����_�?[U�ЄL|�ܷ�����Рd��1C�^�J ��8�(#77��W��1�G�`"H�^os�>������_M}WW!�ӗ�֫���Q��1�Y�gUl9�_=$Z�,�XJ���Bh�>P7hM�$)~JF&=��(���`=���ֈN2��8:8`���_�v�xˁ���]RD�;;;�����bL8ʇ���^�N��[X�����d\�DaC#�:Ϝ����Z_��{t�w���I`u.@f�9J���Q�jk�?G[�܃�»�49]�����­��Nc��FCO�]��I A0�N;i<����KV6k�$��%�.�<���:��==������*��pGx\-�w��G��v�fE�#%2TTb�����7������A1M������ڊ�ܗPE���͈]?�'��B��hg_{ܓ67��V6��/߃\^��� >��zm�D9�̮]Y�3K������?f�f��9Ɠ��-��M~g���_5�l-#� 4���lA��ʸհdc�m2��h��"��ۛ�)�j������z)<�>'��)��K�anD	U�_A�g5�!8W �F	g���'MZM�vy��@���5"���9I�/0�;ux۬�.����A�N�*Ha��46�M��<90�QZ���_��k����y��mv
MoO��t��ׯ�+�˼?R���w7&&���\��}W��2�
�E
�I�Y���zC�Vq8�VO��z:III�+/��v���|y�}�.�2(u�٭[�~:L<�R��%��5����$�&�f d�@}����A�q���~��a"��b߬f�+K�U��S��t"��LU���Ch����2Y����:xP7�op��ܑ����?��k���$~6RH|(v3��7�~��s����0u��8D�T�M�Q=��7����}����ct��is����F�\��h�_xG�u�<07W&+�H 6�ZI9T�V[-��8��kO���"@��(�LN=���C3zCqPgHb�+)1�\�輏����}�>��v��0~ܚK
rzg��%%>�f7*2==�i�N�8\��5���?;M0���Wa�B�_u_M�/Xgm{�^]���<�<���ֻy��綩.�g-��R����oH����? � 4����j�I�l�����8���1����m�\T�q>�gk�01-1[����������z��%(����s^�d}�<=�����8`��XPK)��O�GEP�,�A���/��mis��;���k#=��E/�]lJMO�̮�0��m(�uA��:%���;��I��o=��0Fo����7��������� @�t��Vx�,��g&����<��.d���yVOSRn�Jk))�'�cHS�{�r����u��&[�{=���3WI��.�`D񵋬 p��'']��WM���kyz!n-|��E���^�sJ�X��.%���NP6�h-c�(���$mm�qY���ujj�е�������1f.i �[ix������N���1	�����v�w�c\GO���0̟w�)rߙ���W8�M�������:)�q��- �s ÈL��V�?J[��Ɛ-��蘘��'u�ZxV�1���c�Ų��t���3�e9�J��� ���*k�,���pt���:�
h#,|�v�r�[[3$qq�]��}��\�n����oԋ�pT�A�対��]�f�5A,&"�a`>S�!������x�!��w�uX�&�@vq��5sߠ=v|��� "l��q|_�[�?^�Tt�1fخ��K���Jyh�@$����<
��,|ji}�������F�`�^⯰��w������H�A1tt�+}c?V��Q?��'px7X�5ޕ�h�o��DN2~�8��2%%4��������f�A����i�!(��
u $��SR��tt|�����C�!�Z@/�o+�{�i���hbR&'�(
�e��қ�1�̋\S��$9#J���*�:��P�J�P��\�h��\�2�u�Jaa^lT�.�p�a�� )���f4����W��ǝ�� L���ό�z� ˤM`rI�?o�XWg��}����Ȕ���"��'�3��VT�kZzh�Ǟ�.ZP,�_��U�ЧOd2Y_�C���jh�f���z��!䏆�}�nI������P�#Z{(c���������b0�@�bv{go�8?��~DD�ݾ�Bx�,ϴS]\�_�M7�w)Bk�MV������=>	�����ק���6)�q����o�����v{�Lg'����Xk�
�����?�ne8��M�K�n��Dw&9"�LBK�2Bc1;�ާ���ʐ��3t0ם�B��n@e�**`�RS<�A<o��$�����1����W�I;��V�_�pp�((�ο{�A�w�6B&���ق���V�����*�Бf�]w���♹�0���V��f��jN��:�z��Ʉ�Z��m��l<���_���X�^���ʰ�o�Txl�Vj�-`���xg��ηe��8�����m]�@���6�_����Ԕ>lb���mH�hV[�44���Ԅ�)R�y���L7�܂��(�w�A��bP�T��b[*^dL��+烲��ꊠ���̟\���C�&&W��RdL��Í��0�F��uV]{9 �^V�~~-��E:�
Sz\]N�G3D}�,�jkڬ���Z�?qssu����0{j�(e.N�����a�`�+?���:�R��cN�����g���,~���FQ8�io%G����u9��F8�h9����е��Y�t��qպ
5��c5���S��oߐ�a��J'>�i��Q��jZ{�"&�j,����|�������@g�����K��%����$PZ��lE��Q��O��M�`�(�����11���}��4�V��0�x �s?jC~�E���*�@tԙާJX� Xu�:��=�:���΍��X&���s_nnL�R>�XB�,~�r��Iw-�����O$�6�h�ր��Q��F�皺�)�}�ߟ���������-Q?yr�P���X���51��Мm�u��#ynh�V�Ųk���c͆៌���4���x&��Dz0�G⳰��q��I]]�T��F%� (��N׷Dh�hB��<����h����\

�)OQ�s��������LK�ӣ��p/pL�&�U��V]�m�� ��a�� �S4M�[˓��4��8KT*�4g�U�=��s+&*�Ã-6Z����6mw��(����Oc��n��89y��'$AN��������7q���;��T� #��c����V�/ϟ3�3>h���Ş���#7�{+���_��� ,rjKv�wP8�_jjR��kI���K C���I��z��Z(��wuq�gap��G$-A�I��c���śx���@��׵u��Ζ�^%8)o�K�L��`�z"#O}��Go��)\�li�[�����Y
��Xik��JFn��--7�5����E��pt��]_w�Q�~NT�^)�w�'��؄K�� b��h��j]���͖0���=��Hv9���K6a��k�K����4�j��JKҪ,����eg����s�y�����Ѡ;�ɨ�'�z�i�x����0nϛ��b!�l���-m/�.���D��2CBs'X#�X��;���p�Ç����BIC�9kXY���˝z�M�JI�xQv��D����5�T�[IA�%:���B�l�A�F����A]!�zNR71���R�������z��*M�.O_��Ћ@��im5������h�jg�e
?6f�5�Ɓ�m��������}�$��#�r�Jˎk�]_~����WRD��g{��wvFs���㷁 �|��!mk��/���0Җ��q"��E��G�3�Jx8n�+��_�N�uaH�4��ڕi/�[0�T��&A�S� �0�GR2S�܂bKE�6�t�~=j�%P�90+Kek��tHH��"qyy�.n�K'��YpG�F�b"@ߊ߸y�#��{=�k,�']E�ȴPe���"�������h+�.���"q8�-�7n�fXXZ_��y"mHZ+�����L��vF�5g{�Q)�ʤK67?�%���%(9�i��?/�B������3���А
R��S��)#�����m�^\҅|9�X�{_�P[�ۉӒ��Z|�U5w=�1l|0;����/W�c>؞�-M����7*"n�M��h�T�1�,.r2r��/�X�Ud?*)��P��S��'  ����~��e4ZI�e�������h����sIL�5@1�y�p��6��l�;�K��ixu7���߉t�*,tbz,�D�d/]A�n��&Y��\��\��)G�e��Eʏ�2V��c[�U]�����ڭG-�,(ߺ�D}��,�"�2+�����BMM�x۱͗@oM�		�ٯ`�����-�IK;i25�_����;�(_��u�f�dѵB81u;������p�CY��9jN­wH��1 Z���|Z�O��@�L
��q��x(4����h�p���,"qgU���u ��9��h��~`g?�T[ۜ5�P��< ���/���d�*�u˿C���?��gW����^��q/����\9��HJG�;��ejlx�		0DF2X\�p��Z4�e��
��Ϯ�L�_bT4� �h�$��l9�X�*�B��И�
*�Е�į�8�fnvvН�Cz�-=lI$���dm����{�e��M�
�M#f�k��X��p�z�x/�u.8g�
�����AIO!)��T�č�Zff��y'��܁D'�x⋲���iQZ^u����������sq�	�Ѕ�v|�wr���M0r;�(��}�����z�:K|Hp%k�[� �;q�|�1�>.]\�$4t|תʲַBSh�vXL���b��Ћ���\ˊJ<��
M�ſ-����>��3	ڞϩne&�������i>ܛ$>CfP��d�_��Q���Z@�s�?�����Dc*F�[k�.\�{hx7���u��:�l�+����i0�qK���(���v�3�4W���N�I
�M����]]�=�M��"�`ՙ���b<^�86F���j�*��r�N�Ec^;�����(���Տ]����<�#Ǒ��;���n�&2j��V�5gKc��Á�(̇�[t���T7���2F`.d�/���ė�O�a�	1j��>�L�}s6�mss��F|����i���Q��1r�( >����g��鍉/�'.�;T������2`ND��)�(�eF~(4T��L/?YHIq��p�6Y'W��$�{]���ϯ��`�#G�Ǎx���2�m��!��~�9�r��҆�թ�MFɬ/P�i�����bԨ Uj**�����_u}��ыJ����>F�4{�)9}��P����4����ќ:�����X#�]1�CR�wa�UW�-z;3����|"i@_��DI���Xr��B��U�B��.����;�z�;��A~�ݷK��%i�6���T8�����:X��x�=��4�i��Q?�Bݬ|�>�@��h���֭3ۆ�/�i�ߦ�_�>hR�H��'>�W��XK˛k�ܮ��ZZ����������X�5��2�k�vq�$b�e�"Ū��l��PUG{c��l�k�Cӊ {� ��n�4J(*L�vu;�^�G���Zd�" 8.9x��V���FD�C-���j�C�@&��l��J�M*+5��k�9�i�.�e<�!QQe��;C�h}ԉX^/�E��ep��E)��G~�j�n��j6�����O}̎��San�q����O�$�
(o6#.zz�����bNX��[���M�l�ll�@���s|i|ӑ
E<kKZS�M��ׄ��<36�[�O \�Lf�X�h����_C�_���X&��,��ǒ�.�FƛOa���a�{�OU1/���7�@{x�OSAM�Q��w`�����5�k�AA�J������>!�4�qF7��$� ���t
Ž����)�_�� �܃+k�q�='��R4�kr���	^m��[5�,
�|��3/��#�E��wI8表~��1���.�(�'67���
�}v+#�J��S��Ђ��0��z����T��g	�\��?���{��x;��V@g*��1���`�dC��k3�J���CG�$a�'�Z]�����Eig��P�>JRP~������.��QM���|��fa@��Ȼ>^Y�6����� a�&'�����[���p[��"�Q�7+{�ui�kC�|6袵��Lm1��P�⶗e섆׸Y%��* !_D0���/�oZZ� ��]N���Jq�e�Ǹ�k����Zi��b|���:;-/�O����������]�^����DA��?�V�����d~~q���¢�t;R�-�`��%y����QH���.�qʌ���6�鋵.3EG%^��c���$������O%$,^�1�!
�T"x/ܟ��ΞYT����; '��hJ���#%�8�]@�G�j0��82�+%2��U����h�˴�@>L�lĠ��m�0��T���B�}�6�ݕ��@����ԙ�k���m!r2$��������k��0:L�B�����A&`t��sV���l7 .�_��*��"I�+M���N����&j~��ϫ+CT	V�����F	BN	�@8��S0N��)���<�h?	`��[ b@x�>,����_=���	v�1x��e&���k�}�_Y^�b p�*�g}l����y������,@zl�9p���D�'&�$�&	;�gxه����:��NWAD^��!��wMG�Ga���̇�x2��K��X�f�� "ˣ ii��[�-O�M,pB�e��F+ˋ���Ê
�����P$5��N�v�U:U�['�}ț@��e�����+\Ζ��wL><j��A����tt�A �<��<��6��a#}�۬�3(�-+�ҷ������kkׄ��)�O�lA��NMk&�͓\���L%H��k���=9��u��O]YQH��ڠ��d=�%b�a��r8��(�N2<u�\n��J�{���� ���`W�Mn![:<��^�IlW��w`�'��ޏf�wu�^�g�0�w���(�3:���p�iy07�	��Z5CO+��^C��("�7������DS�:	�Q�Z=n���$l����E0�(lʰ�44����P���-k|�v/ņ��Z��)��Cl���f	�!:-ϒ�}ך�����m��M.�׀vJ���V� �g��������O��I�t��cq��\�fIHI�q�����-I�c�#��4�4v@�_�+*��A'z���fK<�k�a�{.)�N.�0S��1iP������@��<��Z��u"�pӧXX'Z�e���,$�]q�L�Rݥ�V�u��[7[`I�\i}��#��$FF2��\���K�`����N��xp*.*��w7����?}"]�0��X8�+�{�t�<{�,F�t`��l]Mʳ��?��Dm������M�<�
֮h�<��>���_R$G;}<�َ�ш~M'���}���}yAi�,׊FBw�I�̣��e��O
��VL�m��Q�����'-~dS�N��t��uOο
��j���r!�	���t'�7�}N]�GU�����o�7��mnZ�W�����2���3���%���ʭ[��s����L@�h�)��͌��[�>�O^�1�!��AI`�9!��d _�[��V�s��_'ײp`,gc�礯/,�kğ7d�=�%���OC�K�����蕾�$���w��sUnѰ�{�S�)ނ}�x����8j��|�;���a,)�m�m����I)�=1X��N��������%�=�5�<�B'�b𣞫 �*����H�
6l���G����#��8�Y�x��h���9MQ�Q �D'�Q�~R��?�ctW�b^v }	k�9����Çɾ���{J���A'�G������|J�y'w������W�_贮��(h����`g	)(��.���
ߏ�Y[.�v�����	��~4���$%K��ߡ���y�,
�k�/�ΩU��ԍ���-�MA��gB�U ��*���
�Z[�$����*z�	���g��������@d!�s:�9J�Xٛ�����R#�S"@S���E_�n��+��NH\Gt3���z��ʧL��r��q�Qt� zj�u�=�:�&�6|��f�J�֑��(��{��PuM�w�ѯ2�(��8s�W�py��	�$	�ߴ>��Z�b��Ǹ��*@z<*�����rr����x�^7t��<��Q�}�/��)��o����]�q[�7Wl�����Z/{
���F��{��[_J��>  �#�N�%$����C�#��*JI5�/�w�K³���;	��mp~��#H�If�꿠���P���|��4�TUf�'@�T�mI�3|���(��Gu�������4Y��7�����&0H'�n����H�]Mqz��,
���Q�IuQ��@,�C,V�e��W���JȾTT=�b��@� �FQ�};�����Zd������Kqv��-L��$}�w���2V��_���4/{�aRC��xYZ��X�%�q����J�ͳ�!1GM���K�*F��I��;Y���2�i)N"����둯9`�g�݃/-f{�T�}�����hj��U)Wע�JK�lN��ᗾ5m��A�)x+�#[ڏ�����#���5٠'�����_�9Վ3>x����O`()5X^��t�g~E=��s��l��p[�"y��Hk�4������B�]�0R�}$~|L��  ���~�~����4w�)�Xָ=�Va�!�^^��#���}дG`.ɔ0zlu���ǿ('�m���3m����D���f1�7?t�T� ��i/M Q�ꞝu-h� �Z���\�,��a��M����u�8��i�pt���Xt�ũ�J��5�nA~s�:+�_f��!���l��� �Y�I�\���.�,�z�ɪ�����o��d��;2´"�ߌ%P��{���IlR�!���<k:8���XE����4�~!]�g���5��yd�L%�����-��]��w�{��(g��_2�U�e���E����~t�קaa�}Z��/2����v�W�g�Pńw��x�{X��Tw�{�@�U3_%]���$�j���9���_a���\�UAM��ў�!h�O��1�"�C�g��|=�{/	s%O��/�U���������XŤ=�����.���4�4�VR-���h�%� ��+˜�&��;��^�Wx�L>�e��Q�5<vH�fB,] �����;t�a<���P�R�*��z���C�(^��89���8�(B[�	?�C�zY�o
��=/c�"t�?�t�+[����ɲ���>�2��|��I��r��;N��{(}���|м�0yeC����n�%h7�!�dkLn!�%N�Z�	aL��,���EB��Wmu'䒄�Sx��M]>��g�g�NN����� P��������ꊕ���ԏ��H-�����fろL��E�=΍���p'�i�H�VR�������T��'wsN��7���٧�DA��%�������@Cq"��İ�YQ���� �=ݙ�e[�Ԩ�7]ب(ttQ�nH��LJޟu���Xzf�~@0��.��I?Z�}��ӭ!��Β#B����޵�t	�j��Bt��>�W�����Ԓp6�x�8�Z3����7H�\��c.�&J����,�Qh겳׮�D,v���u�O�$�6�����$z����={v��*��א��	h��$�w�f �t��,��_����ٍp�ٟc�K��L��0vp��T�. N+���m�]�{� ���m�'���q�h^�.:��/F�k�!_9�)"�I���H�J��ϟ_2�:l����o� �/^��^i���;1�j�>�=��6�K�Dr�.$0>m���;�	,6��<2;??�Ț�!���׷�͸�o�����;l������x�����㳝#�\ۏ��S�����^��R��>�L�nj��#ܜ�:�?-h-���)a��v&\���K[ŞJ���O���xɀ%�Z��?���cw�X�|�4��O�4�vh:��EUS
�zϵ����
4�{�X����������� @�S�`�)Ǹh&�z�.�����O��Ӝ`�l�FL���i2�Ny���y��F�21��Z{׌��㨕�Ќ�i��˵�ҙ�".���e��E�(�]\��@��+ ��\�T�RxKk�+�#�dZ�+k�<}���p���%)t�)���P��g|��#���	���ieg���O�+�`&�[k�*)�Vgd�k���w��|~OD�w��5��n����5�OP6 N~#���K�(���3���/R���.k�juI"����8Y��.��C�ss�����ș��2�J��	.�a|��;#B��m����B���dL��u<6�wK�z�yHē�*�&��L�����~o=y͕ܸ������x��~�Z`�Pp�o%��V��%�~8�Нm�[4\h-��kp�*�9���ص60�����闱��G8�aDD %�[���Z���(Ι���s>��y��+�.�����(q˯��oEv��d�]��(w/���{��{>��9�+@��tgK�9mX��ɞ�e��ޟ�/�{�O��|v��q��Y�9��nm�\~�{"���)"���|nO>?<��vz�����*�M�z��X�ޏs�݊�ޠ���@��gy��I8Ԥ�*_Z��Nl��y𜻢��g��Hj�(7C��x���&p�b�M�no�i&�Qi[�g@�/��0+8�qh��dٚ70�~~���p��+]����]�>�,	�\++�Rj���Yߞ�c�4���n�����f�8׶H��������Kw�.gYVWq��<2p��3��^v��K<�����|���C0�{$NZ_���$Tq���{I�@����ڬ���%/��@k��&j0�ss����5h5�ݴ��Ao�͹�ϙbQ�Jt��wF\�b��7��DӅ�!��`�R�fg�m���>��+����a፝��̸d����;�a��K>̅V�����ӣ2MT*�{	Y�����Y	��W���@<�cC���[ݎ��V��w�;���9b��
�E�%i��/��s��i�~oRW3�+�[�ML2�w���{���#̖��д���д=ר� �E��NDu�sV���ϪF�)~�_w��>����nH��>:&I@�$FG�UuC|��!J0���@����GS�o.\�鿨�h�Tij��{��F_���+BA���2��}!��U3��2}���_&�^�.:R��;9���i��L ��=;%e}�n�K*�{�ueŝ��΃e�:�ϕ��ؔi���d{{{U�77��@�'��{�B��ZU��Z��T�*iE����B���{Qt�l�]-L\�R?�a��<?�ɾ�b��s>����~`n�2_���-����y�(ߔ���6I�Ͷ"�i�+.qpH���A�!d�U� 1q�ư����qO`ڛ���B�9�z������N���[���/7�+���иDv�!e� �|�x���+�j��_g�̸z�;���xn6�@W��^�@�Add�a�u�"���2⿸n��!�%�c�0����,�]���^�T�I�T�`֏���)�\��@z싈L��6=�-��H�<wmm]�-�����O���x��֖薨��'XAԻ����-��'�s/��<�dC裹g�g�v��'�
Y22/�ڻ�<=�
��J?7�����w~k%O��77�Y��y�S��ŵ|�{��g��9�WQ1@!���}����"7\\�������CsN�CsJ�w�H�&;@v��J��x �1%dc[l�2��g�Nb�&�!��2�#&t���R���V�'�ÎC��v��� �U��Q�Q�뇱�����}N8�����¨(��?�L��J{��dS����F�^�+XbH5S��R��V�H^bJ�Y��/�a\ŧ�l�A�\�w�	�P��z�O�A,�K1����2���F"H4��.�D!�5r��,'�}X~W�ʜ7�r����ωJv�Ƣã��y&�Q��g���ggA��
 ����I6%v=Bpm$h(�~F��"pc��ɧ����VB�=���y�4R�d&#~�"UX�8�ʃ8a�&�T�ʺ}�</x!ax�,��-���@�YTb9�t���U ���;�����r	�^DIADE:E�KP��[)��V��ne�ai�.�����g����8<��33�}�=��y�O�|��,�k'	���P�T���{f���ec�{�ʏHD��*�/��X\��uH�%���ү^���Yȕ;��G�3��R���j�=sPr�B�]�{泛S����
��<+�$�����^���F���O��4�Ź�&C�\1���с����Ξ�O��m+Xl�����(�:��ڝ�GW���.Pvo��yR��p5'��:b�_Y�@O*p��Du��Nt1��"ՙXP���f�'��p�bvy��EF�D�*����w�?����!Z����!�̽�e5�h�z���&T�]���R��ThLR�9�X 7�����l�����NC/nq�i!�u�O,K�K�+�urf��vk81�ʄO־���#�Q��ږ��9�u�0�X�s�]NW�y���U�p���rIx%�b�	�\�B`� �E��ilS���H��Lޤ]<����h)�kf��?���<�e:@��U�紜���u��:�����7ׇ����.	��?^�r������c�G�۳Y�[��Im	j�c�Mv_���k��iV�HP����v����_�:Z�';�����L��=�C�v,�D�`�����`.�PR�h)+IzY#��p���|ՙ/�1`�bl���՞��rX��<
�xJ���וH�r9�@
�9��Z��-�X��6���i��mP���Ik�D}�]�onu��AU�X���^��S`�{R�n��<�澁��R�7a}���~�+a��k��!�v��1*_�vKn�T��>d7���Tn�}sbA,�%yj��T�!�`sݖ.c��nL2t�w`ʢ/�F��#f8,A����n���=j��z(.��v���:�J�͆rqm�V�� R�;6���他�
��Գ�_�����v�N�\
���$�[��h��";���[V]>?�����1�J�N�?��/G�+��2��`��vw�+*":������w8�y2����zh]'�nWex�Ӂ�s�o��"�-A�%�jC���
]�x:D�2ER��^;�Y%������Y�8)w�ʷ w1=�W�������W7�b��`��Wx�b�vw��_����$�V�*�=H���>dp�3n^ǎ��������xNg֍]Ѩ6,��G=��XM�g�|�@R`�&�#�������*|i��%��P1��P:�0�̧�VC8d}_����%w/o.�}��6�\��"h:X=�_B�6�4#H�b��x֡�!��$�p=S�<�QC�А\��>翻 ��R^�sv�A��{��C����c����R;�����Nj�&̐wpwޙ+���o{�5��$�e��:��qK�9o�8�L�'_rC�|?teJ=1R}[�\�QE�f�7?�j9���V���AJ�ȝ�Ro�T`]��D[�uĖ��Ỹ�����(uv�7�'��-�w[Ìg�*��L��A~�L23#p�����ٛ�:�$!#�Q�t���f>�P�ce���:n�R��uH�Ҩi�M#-�)?�_a���3>��r�.����$�н���3�y��F��$p+]Q:E��	�_��6�^h2Y������B��
�f��S�O=��%�v��T�.�����l,�'������M0�͕n�^�&pX���[ ��
�eʿ�`%���ҥxJ3u�֏���+�R�I\�߆2�bѹqDn�܃G��~����S�p��#���jSH��>N .T��+������~��?�U���Zæ�X��HI"`-�?ɐ��XHov��i�"���AoT����UЩĬcUSw�+Y ��q���eN�� )E2R{���ϟ���gu�_��\h~�(��(n/<�:��Q}����� oԕ���^iW�_���)��S���=�>A SR��ʼO�r�0�?���+ʚ��ߺJ��n7�oq <+PU�P�,cN%b,�*��\�8��ܜ!_��l�µ������<��;�l�����c��_���V��y:�$�^�ٟ���`�(?�n����9>9��6����k@A�SjkJKk��\�MsYX&c �&�+�Rb3S����ŭ�}W@�g����R�#�����	4��87��W�8�i�"�.�ꁇ���V�����-U�>XP���/)9c��x���U�:��r/�>�}ZU�v����h�Z���a`��Z��Y卺���c�W����acK��Xp����6�Ԕ����n�H��U�',>��7�nni�i7s)�ھ=pK�Ǯ�x�wdm��~v�}j@y�����cƨ���NsC�껼�D0�sڕ�V���}��b�)�[�L�])�FH2�w����2MȪ��>|W�� h)�h�?ɬ�c�
K׿	S�G�bAA�4�@Vf��.s�^��w��C=O�<t.M����9�-��fG##E�����V��V��-zn5f����MZeE���d������X�]���l�H�+�$|q+�Y�!oS5�GE�yr��x����G�kD/����M��yv{j�uu}�;�&e}R㒦���lf��=\{�g;U2����M*�.ì-�_�%#����u/N���6ܘ��!�	`=��>���?�(rm�j=g� |o�
sq��\@ѨUځ�1|7�����O�]�bN�?�Z���,�T�$a+JQ��{D�Sw�b{Np�D[be������^<�ff�}^wE�_!2�$JKH>V.<���݁�'����� ���0WP<�xo��U�9V�l !��j�VE�����	�:�~JV���a���8s��_�|�tg~f�1%�.�θ\<f��r��B�#�_�`_���*��7F�#JJ"�"?IJ�&��zIAu�Vz`����yHXϔ[�A��ʕ�=���K���hA�"�2$����mO��]V��[�y,����~1Xvp��ZJO���P�I�j�?՛���~���qh0�]�vv�=7u���j��=�T��{:UfffeT}_]�:�HV����:�d��t�>���\A��I��	�xn�6��{��>I:Ï/��i��h��!�����6�#��w!_���8ި��,E��:��'n���
��k��-�3��9%�AJ^��,--��x9�i�1DcՐJ9Y�g�6���콳p����My"����p��v����ڵ�]�R'�E�s�у�3�jχd�/�ʒ	!�㉝jz5$İ��j��E}֟�󊮲3Q�k~�]6X��1�������lyg^hE`vN	�K,S(5�&Z`��p��k�����,Ht�颣��	�%�A�n�ey�\R�����s[��d�7M$/�9���qN��r�}������T�6������5��L��R����&`$�e��GP����И�:�kH�W�v���W���\�°�ܯ��q8-<e�_�"���ú�~_�������ڠ%����S���K������N�����n �������:_1��*�t�_�O��˟a�myn7�\|��@�$ �	
���4��9�Y�������acl�z闱��BC{�):z�_��Z\����șt���W��y�ya� t����#�|���R�4�]�҇^�O��g�ӽ^��`��"�AqK�U�T�຦��M�&��jF��c�}�6�g��u�~{C�'!!�b��?��� S\Hn ���K��]AFy�O{O��13��/x�~y�- d��+��<N�e�O2!Jܕ0�s��S����8�?���W�������~<��n����9c �4�J���q����p�)}���oyi�.�;b6p<���Og�9Z�O	B���>��֓3Ǳ	�
��|{�x�.���J�	��|�>=zqUf�Di��s������y������P�����Bd��nD([��x�)��γsx�R�*����BՍuT�\�^$�O}��"J�0 ��,x*Ͱ�������m������/�MG����cy�M[��J�Q.{+�-t��/ar�[����V+��"��L�e[2��h��
cVr���TY0�D=��Q�3ߚ����M��P�{�:l\ 7u$�V�����~70��Gs�W4o=qj���y����7����f�����1b��D���XTbd�T˩��Y0�[\��tB����C/�`��)�_�'0��d1%���I� �y�|��ı�EX�,�+��H�vu�=�7�rƑ�ii��y9Q5N�s���:�v�L�n ��7����4�f��(CƧ����v��i?�#�����Iۅ[(��9^[�_<� �{p��2�v�d�{��|�)�)����1��$Q�2rEV����@�C^G˷,\��]y(��m�����,�Wb�����w��ff^C�C�Fs�2d�F�
^$�\�++�Zδ<2@]����\2��0��¨+�Pj����F#4������*�ǃT���P1M5��>��eQwF#�]�P`��w0\�̬�&Es �O�������.��*j[p����������D�l�l5���R������4�D�ܲ�Ng�t`����/����<����ꥊ��;,D��������!J>�4����}�s�r�����l�;o2�MM�JA�ƉWe>O�H����-�1]���j�k�[3�ƽOGmq�#օ�2��+����ػ��СV�d"�������$O��@���V9�0 ;B�11	�f����ZWG��LE`a)��1�(}|܇����C��o�뫬���Q�p�/X� )��n�\�(Ri��:�=����f�~-�	�[j�Se�$��{WY�����ʻ�������z�v��`e���m7ƿڵ�.vx=�1L�r��@����vK�z$c!]*\�ݸ�j���щ."�ә�%�d�EQ�c���\n�W���j7$0�'$�~r�E�N**E����?aT?{�ۖ�,=ѝ+���ji���]?'������L���~��m�e0�����:�������� ͆����}'!]%:rM@�8j?R>����m$��~��4T�`�f����촄_�Y&�jj0�r�s��)UB�'5UKk>��iT/Z��>��1G�%Zq������!7~Y*dr�v<�%�	��O�wR�6�}��t,3��H��ٵ��УNH�zc�1��~�-30��[K����D�K�Y����c�)�Ƴ��iN�t\�&��B��K:(��������M�|,�_��3MDw?WK?�r>	�l�[�|h3mtL���v7�rѱ��0J�'7�hՌ���yd��2��[�}��*>���?Cg�Fg��{	
��Xo�#"��AR<�/7W*������j��� �3�)�~j�<X����)st��}��?O��N�Q{���`pi"����@M���/���آ��r+y�� �'n88��8������{tq�Q�L��`@�q��w>vf1wµSR������i�́��^����+1 !����U�k2J�V��� ����F�
�Ry�;Y�O11��v�_p%̿��*b\�;��A2KlSIme��6�������V�"�����+6��u�ȫ�Ulum0�'ǽ"��SS�~��)�r1�U�K~qd�˺���i��P=;Zp�x'&
~u�n���&|�
����QYw��7?�bLZ�[���Z��k�U���ANU���7?uV�t�?׾�؛�\U��£�Bub0}5������{Չ17W#�$��ibl�(���h7���1+�ۈ Z������c���?0�;!��6<�uu� ���Ɛ�GH����&��B�1ܟ�S���|�i˪v�x��6����	��dn軉sS��0�N�}�ÅI�,�,���b����i�!���� =�l�g
`�|ߋ���'���N+=ۋ�%�M�0(�M8m��4+�g�!%���N����i)7��Bk�h�W�n7�����jq�����+$�1��hL�����K}� �eU�!�Rp��6i(h����_��s��
t"2(J��������C�z��Ps�߰+}�wAJ'h16v<�n��Qا+�2�b��s����_���?sD�$dO���M�ڝ1����b�R�s�ׇ�%�.³Aj���W����X���V�7���#��]ó�h1팒s���x��W�\��8���pMM�ט�@ʄ���'��F��!��=X�@W#�\*�[z�iC��{��4�I���?b:�w�/n�!eE9��{����3����E�b�H��`-�+[^��Aly���չ�Fͱ�>�YJ-���(��F%��/:�dp��>�/ ��x+C�^i	���q]I"�9�B@?,�b�{����Xl���h���B���i�;b&����Y�J(+t�!����Q��J�Lzv%����Q��F ��]���$;(BO�Ř�q���yJ���FY~ ��T��s6�â��o�i7�f@~<[���c�>fwu�5��`�
��7�$���%;32*��DCuL^Du!Q�y�C*��W����P�E$����W[@�H�G(o��~����������	L���P0��b`��tH���]NG*ͨ)�^ڌ�����jH�A��z^�xu��&�aK������#�Q���Kx(�	k���x�u���T]'�v=��Z��=�DH2�����ю!��\6�}�Y��gDM��,�5^_w儾���d*�ۡ71��[���F�+��>��2��1z�V�.�'�t�2���,YԵ��BT�ʾ���f�?;Y]�^�-6]��p�'��Ƶ*8}T�����݄ZqSdi'N� Fql�i^��::Fʑ�}��t�{w����եW-�������nNz����G׀Y�,/+�n��e4�!?�eB]���Gi��4-��e�����3�~}�!��R����MM˂Yh�δOmIr�����-'1��
'��>��9�n��$nnjcMҿ�,�1:�
E�Ʀ�g���)r�\�����ec�j��n
((*�]���ϳ����G���9��,/�����j�t�j�rt������ͬ!�؊P��6�`G�gᣓ�P��Ĵ�y�'A��G(uqޖ���V��%9�2]�=��k��bu�5A�{H�]gwp������7�!#Tw�m;]<�� #D�Y�tB`J�6y�ܟx*.frd�Re���j֑޼6�]1}��3b��C��(/��ܼ�i���>їH�|$��yfq|�'��M�.��,�_fNM���?"$6R}
��9.��@\��=?����2�Fs;Pmj�023H�tv��`�}�������=���Ѽ�#�d��
2��ݾǏ�����?�M��s�!��bFjB�\��O�J�r�񣝣	�TDLfU	 R�r;I	]��t��F����_��n43#pp���<ݛ��BÅ���s�0	�\h�����~�L�LKН�^9y���'�gw���O�6� ��P�=��!Y���
t��9 #�}��s6G-�硰(&^ݫ|��{�sQ;�??�iv��귯��jT�{�����d�ٴ� 3������*�,������)C��kdEG��2$0:Y��\Kh}�a�3���5e�u<\�}�-�#%��)�1���M���Ѩ)ٛ%��"�Aj�~�0����۾�K�ٺ FH!}�`T�����T���L�9�G��|㪛��Bc��EF���|�I�\9����Go'O/;?u�7��>�#����� �D�������"G�B\X��:UK�����DU���_G�n5 �%��SqJ9�tb_ϙ?�����j���u�yX���gCE���M�:�;ɫK҆�ӹp�`��Ų�.��zL�? `�E��~�]���}�g��L7�i���JO'V�ȟ�-�L��h$rKCS��2kԡ�=d0���A����ht�J3j�~<��}�^Q��6�РP��yy����du:��BQ�">q�c%��Sn�t3�n
�@����Ё�z�T�""G
���dyu��I�:�Zna��c�a�b��I�2R�g�Ǩb��\\�ڳ���kS+�1٣���(��.�H����b�v����>u��ϝf���7Ǥ�p�<�BG!���M<�vO��NIɰ<mi��8����}�������W>�u��#3k!��3
�MZ�΀����8���<�a�Td��r 쭿uBr�!��奬�X�m����&�z�����&j�8����A����Ŗ���ezŬZ�}J�twG)����D���ҐŲ� �u+������̼������w%��| �b�	2<s:��D e���p
��5eܘ����!Jƕ�w���͗�>�U@��o��/4A�o2n�|y���P�6����0�z�����8�EeQx�P<1��~����[�g��b����a9�$j�n�ru-��=y��=��5Zu!�	7ξ�7�i��c���!DI�2�X�K�!�][s��w9ZT�(�ى�|�N#"/�2@�a�����P�Ú�Q+��it8Q��;R�#WN��Z�'�)� �	��B^M��O�vg�nIJ�h�Ҏ��#�	�7�]��?�q˚��q�5�!::��I��%srl}�����5h��0h���"���us@�*]"J�si�n��n�oM����u`
Sj'���f�~��h�q+��i�ٹ��l<�X,G�����u=��Jz��1���p��Rɏe#r�f��6��C���I�de=�v�2��U�E�������8�>�@0�-�b4Szo����Z���M0���_�Y4���ai47/M��T�cb���{o��#��D��guL�rۉ�YBDީ E�!P!'.�O�u�^�XLy*`x{R���?:��ۼ��7���1)RP��|(J_��Д[�kux�����tEEE���c@�<>�V2�+H��r����S�����ǒ�W�>�	_v3����+s�Ю�ANŝ眸a�)p*��H.v ���1�I���En�3�
�I������Oo�b�t�u<��\rW����0��V&����pd���[�ۨ��eSa��I��mU|�N7��!D��S��D�ff�,|]:P-� �ws�CR��lT���M��p���u���}��U��ڋ���3��D�������bP09M'Q�V�`�.~͆��'ׅ���B���^�U��(�8�}�3/�n�ʿ�!_Y��:����P�<��W�^��z����7�4���p�GU����	uvu�H=�H=��zbS���$ڶ�:7�é�Ԭ���آ�_�=���1n0ra��d4��z��F�"!.h�I�Χ������6�F݉�.vZ��<-B�{��'�Į���&;0��YoX��n��){��Jt���g�H;�W��@m�<m�R=8OS[�\Z�ȵ�,��j�g�c�O)�1ZS%7�+�>Q�˂p���ӳfoH����AA�xL�<,�m���.�B^�i��1ϒs��kOy�<�!._~8-����-gv���=u=L�~{i)�q)��F�����gVK��K~w�ܷӥ�-3������7�R���E~@~��g�y��N۾���B���<b6��,"�bk�'�C3�B�AY:>�#��w�Q�و�P�B�_4��qX?c7ư�)o��U|���|	��o���V�Z2�h<�?���U�D��o�va��?y�7P��_����W�x�^���q�װ� �:�֬��u��Nb&D��|�%�]�r�oENR9;��ȏ��߹�8�������1�,���	�{�oLy��|���Eb�Ϋn��%f'Sm�*O~_%���^DYu��Xy�)XHz���Aj~�(�h�q����~����0�v����2<xx|T���,!��)1�g�w\�L�G_G��`"`��[���*��h<"l�2j��pГ"=nNBt��>���SX>ɘQ.�U��HR������ގ�l���M��n����uԄ�b�� d�z��Sox�[~p=��*�0��z g��K�����/Ưr֐�_��a��_�)B	�-|�tq���i�����W��Xd[�Gw?���6*h�z��x4�(�݉g[���=duGr*U�?V�6>6�L�ݒ�����_ۣa���	X��n����V�̊R��l�5�+.c⿜6@�����ƙ��;��yC�^�-x��VC��WI�n˹��5%�\8E�V�?K=.��埏��>���$�� �ԛ������r�o�u[q5����O?���DM~�8�۴���=Q�,�u�$�{��H�i�:�9�����Tkn+�B�D:S��ϖ�ͺ�5
z>�W�E|���^�H�VK���1VFRϛQ]�*���-C�PX�^s�����B�t���iːV���;7^�6Dbt����/����#�Z*)b(�(�!H&nn.P��w�×�x����xSS�`�%�RS���I��P��оJ;���2��c�������E�+-���P֨��0�e�1�r��̮�^q��Œ{���_^���\;o�5����4�
rΈD�^<�j�V���[`�����җ鍍|u�t(�P���C�$g��q�k�qQ�)�`���G[��[��B�M^�Pp�DFy�{�����>�0�E������z�gޯL\���2�V˪���x���NK����S EQq����$�[<[X�m��tk�a6j,G�����S���b9Y\Ћ&�:��;kW�d5�;}��#%��,M��mr���11C����7[�/X/w���G���O��]�u�GX���W��:땓%��-��;9O�yAZ��#ڠ�@���8 ���q����Q�rλ�O8��Ū�v�+�2'�&u�pQ?�2]G�4%�*���>u_h�a�k��p�Ͱng,�5Lo>��x���ShS����;�D�l%�؉g�)o"��*횳G;��_cM٦qJ��mp;�	A����}KLO�m/�����3�*79�
�jN�q�e����e���mw��	 ��ef϶����p�׬wd-��C�����Nl<�Ȥ[����� �"N��	.G�pt��%şf���)H��ĸ�"7W`Q -�C.vH����q@]�x�jd�!��� s��9Z��F�پ�Q;Q�W�Q�̋���3h�5XcY�`ڝ�MA���Dc��dl�^���*����"�A;���iFT�G����N�]Y��)�Q9,�4�����4>�y��g�on�vN\��C2sN���"��$����������J�j&Hm+7�L(I\)_t�}(Ğ�Xf��T��j�UW�o�9��S������GGY��r�ŝK�5c+G���'-�J��J^���}�J�i��Li��!K6.�����T@Hb�#�K-�)�~68(s����6B�F˼�UJ.s�V��[�Y�B�N9Yd|���<��Ȭ�#F��{���qv ����"�dGs�0���>���i	'.xo75���aA�ؠ������v{�岽I���M�%7��iT�9�}�snX�h�7(���ѵꝦ�	ӿ��{$cŔˋ���r�����I�U!�mc�
�G��A,�?zR�/_����@�#z�^e�."�n��i:LG�����A�a�����\�{+'���?��nZo��VI��9Y,B7���@EG���v@P?"��Ŵz`��J#�T@��~-WįE�H�9����F�m��Z�R�����J7^����;"r��A���.R�@	�C�1ж����mm�\X�g΁��,q���-»\��/M�
�F�����9i���$���x��ML�(<�k�dC[n^6�Y�~���t���9CT�T��:�V6҆&(mdt� ���m���!�G���4�%8�� ��̓�?�V/+6����Z	�o����w;�[;ItݖB��aPQV�-AI���� �����n5�s>�^9��.��5��@+�,�L���Ifo�b�j��ˌ���+�����OI��;Vbb�]�q����K:&S��Ϲ;0u��3��-d%}��E���� � ʶ�yq�'#)�f4���  ��θ���,�����֋�P'��Q�v���"��KpqB#e���14T����̴��#�5��*�Pv�����i��a�a� ��gb�
�\��S�o�1���� ���w���m�iv�Y$K��&-�;b�</��fВ�R�d�p���o�o�b��E�>r��4PY�L�#�g����S�z�?{X8^��B�[�Q4��TZ    �֕�7�������G9!(�(���ZP��G�a�+^����r੿6�9�O��V���n�
��K����dBU>*���s���9Y|��!�)|4�AbΒ�1���j����w1�7��r�-pO,��7�+���ȣ��[	@��'o����fB�ŕ��x�I,��� �u�nA����DS�`%P�
9���x��d��ø*s��.���V���YɃ�)�E���{�E�JY���*�||'��N��R����"�;��YG�l<�Rt��mHS9g�^�,�a��b`���=\���ѯ�tB�w�O��Khh��~L��uy���� �,ʉ�JYq��
�y��m_�~��v�]OĎ��������� h���娼�ҁ��J�6�
�(��&����`*��<ˏ���LJ�-���{8�h����i�T��M�9�F/����Ncz�k&�b� 1I����y ki,-�p������x��L�@_xT�<���>�pM#rif��m�,�lǂ�����~���:.�YϺ#�� ���]kF𣰐�**��Q�Z��vʼ���u�D����^��n�����b�y�d���M�l�Ҩ^-�w�e�(�x~���pg���Y�G�8[3_���]��`���Nօ�>L��Hgݮ�p��Ąہ-����әRͮ��T�p� 2�:��P�Q�/3���~T�߰��^E#����<��@h�dQ�ו����	|uhzx��<��r�w?K���'O�Δ;w���~��!G�����uU0���?m,���(,?Q[
dܷ���qӖ nTt�<?�$о?V���(��P]9{}ܬ������נ���N�.�\Ov���Ǿs3\��ڸ�~ �iA�1�G����X�I��&��A�m�ϡ��-��Lq%�i�+��3e=NFI�*V�Y�7�O<9"�ac���1�L�)w�M^&�.eX �Дկ����j�����DD�SO`D5������%`��Q�j�I?����`�$��`�� �n�wet�����(��K[7<���n_11��!�%}��b3�PGqӏM�[h?�ɐU�[����b�15^\�u0J�U�V�����}�yA���	�K
Uj�>W�;K� U�܆�-�'�x%@׉HOײ�U�8��jm�8�[gLdt�h9='!���]!�P��]U6��H��j�f+�JLǛV���U��8�:�1�M�4%t��%t-<�;m�t��h*�|��=(�K�'���i*Aǌ�8�EF�;��� �8܀%�&�Wr�L~~�V!��R�B%2Q/r��dnC�k@�U�RwWב�󍍘`�sT����Q�o��,�����\��w�,&Q��Ѷ��Ƹ��&6B91����P���<t�y^���uT'����0���4��p��i���`Z̔9 \V��9Pԯ���6޴T�<ݖ'l��$��d��2��RS.��E�1��)B�7�#캊�7/`]~ ;A�Y� v	��Dpo�����*Ɔ�8g�����M��n?r?��,A}!MTaM�h�MEN5E�*��<���hV���.���婤�蓒
��?�+��1m���N���h|*W�Vjl��ԝ��;�@�/$D�F��%��=��)�I[PR��!!��66�>��;�MB����o�Pw�4>^�ML�ء`E�����v��ˑ���x�n��Z��8��혤Z����m7�=_��p�׻��{��iۣS&��%0����Z��c��){�-:��D�@�a��^��	]!���3-�6!xO#��7�.8O�Wn�eVH��j+	A%e�~� �b;Y�J�
��a!
�GǕR�������#L�y��q�`���N�~�')�� <+����_7sd��Ɍ8��� ����Ӧ%� �復�zV`qf?n�M9&H��j\H�B��MUC�5bl���eծSS�v�UӃ�^�-��nωUx��k�N���^6�UT�T���u�
h��x��ǃ��.�>$�yV� �0�_�ʷ��̧}�4O���D9Q�va�>Ww>:Pр6���O�n#�hq�Q�>�׊��jV�@آQ�Ɂ6ѫ��b�����'(rNǯ����]:AP�Ol�ٚ��h��!Ѫ��:L�P.S�I:�O-Nt��-a#5��!��M@�N;#-��=��P�O���#�ӌ
_�ĸ���#�O�n�X���;GXnj55��8����~��U���^?w����B��w��	�л�� ����Q�Z�'n{ykG"�f�k��Ō]�R����vp<̂�=��=ᆛX��/�X~�L7Y�}e�c��ƈ"��
v�5K��ը*�q:ݒ_H5/�h�(�98,�����
`�ffIHjoy"E��<=O��s{�R��H���vff.\�����ꏖ��_�^���a���0\Z�R�7�"p��Ӄ��y��-���I&T���<}@Vs����n�[��c�C@�h���Dv�=q?[q@���PVn�p�,�V=�'x����x�۠������9���V�����9�'�Ϲ���Cm�ﾜ0gq !���[��kk?D��(@�·V�D���������_r;���%�"	�I�D�ftT푪��kh���5V���-�vz��R[ʏf�29 ���G�P-�=�'g�&������2�Dk�O62V�$o��3d��O���4�߮�h5��U��dz�;Ob��g�
0�F&�Gp�	�r��Be��"���m�
�67'���':�-��;�?�D;������5XOԶ=��Y�F�^�tE���������À����h����7�٠Ɏ���Ɇz����2�(m17����C�n���[.w&1�k�f�Mh�.X�f���1ݿ��eh�Ȇ1�jn{o�e_�Pff�����6*BK'y=�97�%pO��HV?�m���A�����S�bo��{��Y=���aݝ�"V�������E�EdJJ���JS'w�_{\�?�S��K�c@�YO�RG����N�"���2�+��%���������nO��*��0�Q8n#ë����}d����@��N�TI���߀՛�&]�d#�@�9:E\�J<�k��P�r���SV)l?�t�J�����i�`#��^g窜�d���s,1gϸ�����wn��(�Q	֑-�tq��B���`ny;	�����G�kif#�A�������|�v��Y<qόi��hW�d�����n9�����T�ҥ�����c?Rz�VJ��C��:�Z:*�8�>p�h������������:Z����Y�9/y�qt}N��#)\�I���sA��+C���M�/��1�8��ݜ:����8� ���KCh{��.	��mN�ڿ�ԓȫ�r �JK:R�g�&�E�J����jg��	����n��|<;�V�M�j��ng���@_H�huc�)�Ӷ�\���OZJL-{g'$ViS�u��s��[���(qH�~��a/�BQ�$a�m�2���?�T��4��~j�B*�N�w�� ��|��OB44�TW�W���FrwӀ�z�`��=�G���vT��{�m��X�Y�v ��������E���0��1�`\����ЕA�ٿ���Y�sw���ym���I;x�c9�&�(���z8�g�_��=�2��o�
mJ���P��/c�o�gM���?��������[j��ں�J�S��i�aRTp��$��(�d�U}�ͱ�i�M�٪$H� :M/��9YO��MOM!EV+��>W4э�늛:;)�.����^�����#��z�2�����i��}�����F՞f�2�6<|�I�FJ�E0D�]q]����o��Y/ʁ�EU�6�"GZ�F:�C�e���_����ڭ���2�+b0/��t@���E��'JF~�����(�>��5���a�Ձ����ۀ��r�!C�w�����Do>���B�Ѿ�v�T�S�]荷K���$��D{B��x��UGG�rSu=ozb��������3?��*�9qvؗ�Ϭ�� �`h-o����Y@����d�
w5�B#�;���PPgS�ө7��?�r�r{d�[��,��Yq�����9k�C_�#8�3
�裣���Y8\u�p�9B\��{���}SS�B��(S+��ՄAդ�Rn^�\^Q!`�����y�%`o��Ȁ��H��<_��z�j�!����R�� ��8EޫJK�}���{��v{�_������H�F-����l���5,`nn�d�G�/iU�_YS��f�n|	�G��rҿ�^T�'�z��4��U��L-rh/���R��ɉۣ5�5�9!@2�w9 �c�e�Σ[�b&ȹ����˝��3�s/��#��?f��������r���j��y�HL귒E�[0����e���K����e,T{F��H����Clz:�Y:�'}A�L��\���ѷ�>t�P'�������xyaGiE0=��97 �z>R��{�V����1v[��CDŅY�j�$��Y��q�`���2྘����	�k��@G�ch�ur��0a=P���%�a���o��<�r���60�uKb""��g2"������|ǃ���\�DK��N���7�@IU�1��A�r�w��E}Q����C�:�_��n{�v`��kJµv:O[3wmD1���u��F���s��d��g�?��t�]���$i�z��*0 A�<f��_u�Iw��+M*���3��*�KF}�ſK;�Gr:���h:'A祬�lH?/;�.W�.����c�nC��C����K#&�e�`e�2x�᭭$�����^����G� ��j�9�}D�,�M����P�"���"9@�T�O�Z�r2g	�����BET��ɮ����9�A����
��R֨��rҧ���-��o�im}IB�ݷa����S�d|N�U�d��F}�J���
��g��qڬ&��3= u� ���d�0Q[+��W!��2Ն����F����0eӂOrkf�ڱM����7*���xLi?$d�g8+���,��+���-��Q6�ͺ-�����I�ˏ݄ޗ��v�V�	.o������ݐ"`,Ks�$���Vƍc�` �́�c6Z��TbteU����5�޴��c���N�m۫<xv�qa	q�g�1܅���������2�uع0t�d��{9d��FI�p���t��0��u}7j�nS�<�M��������7�R�T���b7��ka�ग��ww�rV^Q�`�:�N�Œ܏�Ry��n:�y�+����FDཱྀ����x��R;��b�۵��e���ߢD%գ�;~~���0c��5,�f>�����I��p�����̇�`u:TN�BB�����P*͌���5��������mZ�8��V�d8�aC_s��`z�������eIvܰ���R�qF�Js���j�VHJ�+��jಉ{�5.΅��g�/T�0��H9��.����;��<�����04+"�T�l�+H���t��1�(E��t� M�
H����A��������K�<1yvޙ{��;3��)�C�%��<E�e#'�8���8aR�%��p�&��rF+:n ��u2�תk��z�<Y8G�zEEm׉�;1��(�9)��i���X����G���=E"�\��]�UK�'�l��.޴�7(��9�88XCB"��k�s�K��Y�i���<*Y.m��C�� �x"y0}���Z����Pob�{K��{J
���p���#t9�@b5g�Ͳ��7$��%��r�~���<�II1,�8 "F�#��ĭ�<O�hm�w����\Ά2쭞��sl	���A /�.����S-Ʊ�yĚp��o���x�F��FZ>�e#�(�N���D��@A�2^��%6�oLbk��W15�]@76��)�����ߛ`�}�8I�{waJEzv�KM\X��y8�PSC�|�����������"��{�ap�M!Rh{}��cK�*zyܯ`��`�6l�=��h����V���O��4T�KW��S[Uz�}0���Z�Ͷ��F��\����g���Ȉ��9O�S�V;���BMήG�Y͗
�b\�����B�l��)���.e���	�d�~0���W�+����?�c�]��f�>4�u".��l��/����D��Esө�c��BY{|�n� ~I���V��N�nQY��6M&&�����C�~��8��i��Z���Ы36�t7�tnY@5����m
<���F_4�w\�捖t zN� ԕ%���{x�ۦF������Fb�M�� �<�=�%v�KRH�v����$K0��P����|5: ����	�"Jn�}�ίB�Vo�%�D�FF4�͓&;��c��b�a���v�${�$�X�g��E$���� �Vz�������_�NQ�����ݜ�W&����eNY���Ձ��ӺD�C��($c(A���e���3*��Rw��W��;!��b��2-ҷa�4{�xX%�$����Z�Dj�f~����V���䎼�~��|�R�����+x꠼�J���%��CM��~|۲�5O���๞�����ɹ�8�7�w�V�6�9ρP��уM���cK*@b�\�޶i�FX���������e!h��G��g �а���΋�~����\�t�wYF?2]�n �Cw�� ������Nܡ�BAT��è��1i��k?��B�4�`[��W�S�VX��ş?�DϽ2޽��w�����%��|,2j���w�7A�4���S�.���i0q@�忴��ʋ3����n�������U~�y��rR�?�u�<��tK86�\́�� �ŠF�qG�/�q���Iڻ�Ѫ������b�pY
�i���,MH�����X�Ngv�::8�Ļ>�h#Z�c(`Svt�ԥ��͗rv �Y9����1�-:6�+�Ӝ�֢�Uz?����0ޟ��Y2�K/�;.�=&�.JJ�Q+�#���r��hW�:*\ĉP���nu|R��=��=�cc���o�'�J�?w!{o��H�YG`U���R����镏?�����;̨���g���z�6B�6t�3$��A��H���zA3 �9O�C�.��ď�њ����ƭ�p���}�^�w�ѣ��	7���~�Ue��BM�:�7q�8�M_P�C�(���z��_1�� �˾�����'G'wCf3ʤ�F:Kڒ�E�![�����әz����W��Jf�أl4ZAbS�4m��)�[����/~{m�,t1԰��DD,��� U��7lGߊI�Ӳ��~�	$�ݸ�b����B�L�q���É�)�$W<}�i�����	�������"�b�g,��Jk˝�A�"�BBaP���q��~�x�4ָl�������Uh��SK�N+�<�m�r�P:,���J��ԫ������O�o��DD�c��Z�g)ҍ�I��޾�I��g�n�l��r{zvFYY#D4��l�ф�k�%cÊ�S�XB���%�n��DKn/�I_9
�+Nc�i��79�v}�bB�ϲ�l��m��`x;hy����T(��~�$�c1��Wc���S<W7;&�s΁Mk�Ub�L}7NL0�	��(}\nQЅ=�LK�$ߌ����c���,�\Jܖꇬҿ/�EF}�q9���i[93[�~�mj:�{PԱ�d'7v�
O��1}�TDa���HQ��F3xz�kwg�����&�R5y���$%Y��D��(����R���y�E���뫿�.�hu���Yƈh���c4����Z�����߅�� Q�,�8�hП��� ,r�5~{�:!�-�����}�+��K﷋����GY��E�{�,�P�r�Z�µv�ŋ��ب�^|k�����!���{B�r�7~��a6 �}u��Wbj���2'��vᑟ���i#����ST�X�"b���~Sîo�tC��X�������jf}�lM��a�E_p4Ɇ���y��Ҵ?�N(Ei��U��B_Q�Oo��5�.0?��W236P9�C>�x���.�_�ca�Eu�67�i����Q�xz슼:�|�v�7�_��
�Ѷ�[�|��xVԞ;��^H�w���C���Ӿ6e1[m�0�g�s�P���M��4�1���`���ˁ{��l�ҋ	� �� vP^��	��aߠA��K��}���8�8�Gܹ$�^rcB��2�N�� f�u���%h>���EW�a�i׋4p����Y�G��^�Ǯf-�T��������}y=�,�*eVQҟ`ө���q�$���q�w����@�����Bm�
�l]����d�%n����s�COA�����8Q����x�=<�u�����\'��.�	�JI���z�$�t4�5Q�_p��!�=K�|���W=v�K�±� ��cg!�]�~��AA�����B���6�y�V���w8(�Z(��V6�额v��ފϵK���K�Y�|�1Rػ��ߎP��r��&��P��<����갈E��[�t�wD����I�;�jF���yc/Q��`+K+2�h��\
��.���r�:�`��Zb�X���ŚTib��xgB
`�v[VA+t����]������@��$*��ǆ� ��#��.��.��準}�M�!hEޒL�3"q[�v���e�G?�D��on4A��V2�(�qlY�c�(��H�L�,��]\�֬���i��¤z������4ɫ5T�&��wYD���:�z��O�W�l��>�P���W���w�S�I�NPV�����p�)tDu%+��!�}�F���l����9����:�C_�p���Z����z.��n�J+c��ӈ����K���y�h��
�'6�}g����@f��������=9�K�Iv'�$L��e������]�s��SB�y��v�E\�7�B��wJ�}b���E$�4"i鸳�O�r�������Ob�:P�����B��v:��K�	��@��7�=>�m(�&�a���6@E�r�E�c`��U��������E�ӯ��h�B�ÍEZIc��RwG�s�S�En���$]�tjrD�n��Ŷ����=cά U_tɌ���&@�b88  q���Y�F08���1�[ �x|����x�;�-qb���'���us�Sn����q܉u�n�!dkϰq�~��e@�hlh���Ǣ_�l�!:�㝇�����K�8%o�x
@�����}~nl�!��L���'
���5x�����|a{SY��2��gP���x	vdа�	w��#�IJ������ P�`	�-ЗM�|�����	�|�އ�a�e���u����c/V�b�ޙ)v=X����s�oEm�6���H��]���aUA�	��l@V�h��o�$�l�/���^_�����b�+�;��aE�oT�B��zI�<7N��йW���.��Ad��V�i���ǋ�	2mHY3��g�+Z������
�3�,�;��I�d��N�L�b��j{��
�y�ڤ�^w""6b�������;=�e짤Y����*gAڙ/���9��J�d�
�ׇ��7{b�ݺ��,m�1�Qo�8��3$��g}5?�H���WRc�G�ñ�i�{�(�-�[��������o�h�q�����[F)��H�[����|�p�������E]�^f8���+t���M���,9�H�[�0���twgĝH��-F�j{"�w��B������1��� '��I�c��(��;eq\��zn슈�d߾�~�;߃?�z�J�=I�'�I�[u����F�XП�9��\Bͩ���g�T�ywR:���\t�K|}����j�7���[i_�/ǿ9_^��~��(U�߳�,ӉKK�Gq0���b]�~�u����:��k�]9#��P��Y�������W��}T��y�:)K�rDq����܊�I�pɩ)C��/�6�N��a����5��m���}�����(K��ݑ1H�1�����1���(Ov��f�!{��N'zZZ�o�^��l��N~�f�:�%�V���B��VL�J.瞇Ǜ��vvq�g*��abd�	"�����������/0)c�����Nn� �8��muu���J��׆�U��h}��W~׍�.;�z)���\����\�f^��4�;{C����;�X�C��xx��g���k�՚[+��{�k�n�̺!V6�T`��n�f����;�\��.��Ǝ9��^֙�n�*��h���k�:��Yп`=g�Mu?��I2�d9,'�z���/���3H�����#�Ǚ��E%( 
�ru�s�%6v4OsZ�/g���۳5��s+���[�Lj�}�kS,��dh?���&Ox��;�I�����ۛ����[[z����AR&t�_ъ7ܰ�H����/�t��%f��l����Y �/`E��9�}�DO����
�s�4�W��g"+���;�j��>p��
6���ٕ()��~��m��{E̋��y˓����V=�է�O HF>t��k7VBkC����|��lt$: �����⢞5=�^o��3��s�Sw����hh�Q��`D�~����C%R�O�I��SzI����/�wϊ�UQ=�?��c'+�$1�U]=����,��ie��L�E�E6g�To���4�ܲN+��%g���f�x���jT��-!��ِ�	a��C@b�m]~��4d���؝���[�f�㑕�X����>���a�m�S�Z�f惆��U�"8/8��s�	m�<���j�}���W/��m*z�.���{t��H�-A%;vT>��JxR2��;`�귳	ņ�ev�~�	�q~_���oB����Q�3�x��c���'���*]���#��s��I=��e��\�H��z�t�D�{`��qq5!���ƛ��[[�7���}1�ЦT_qZ�d�![ ���!:�F:�M=
�r�D���ya��{����b>p֤dۑl��#�
�K.����=f��*˗"l��j��LG�:Q(�V4��^i�S��s���j�
 <��rH|�r�y�
S��9�)G7��[I�81.���\�r���'��tXa�23��c���dLA��s ��@����_������X��P��CF������b�B��)�az�J"���ޮ]#�{�����)�Jzazz�;ү���1����e6zU���b����i�&��ГD ��I���,	�.$�=�-���tR��q��{=qU,H?|�1buu��S#�T�;����R1L���g���]�Nv �Z��]���;3P�.]:�>1��nn��Y�Ei�fxlF�������glc���:2`����hii9mp����?.FŒ�O�f�LHg�L���Q��<�J@��T�\���V�(��q��������8�
Б'n-��e�@��<�ttTQ<�~un�� ��\��f�O��.;�0 �^��YR��[/����BE��@>(�����!?�ʙ�X���`2p���LN]��-��R��d{JiΥ%�j�T�eS��[Kg��<�cI����gYE�ͱ�Gy	J�(���c�r������g�q�P6X�)�֎���W�e�o��2���'���
�h!�t{ʷ[�����ji)�|��D_p��2RZQ�ޖ����K�����1��s�Ʊ�_<Y0^;�B��rF�Ui<�.h9ʶvׁ�O �z[��H�ue�������@!Ʊ
��������t�����LT���U(,�b�l�uZ� Ӳ��'��S��D���e�Y�by=T�ʆ}M��7L�P���^�D�d7y�CK�7�-tL�s������*�p'������;�&�=�_p���%&g�z�]��HG�Ի�"��O=����E7<�쌉 R8�<�xWZ�;�S1��Y6;o�L/���^���+�4<�|O��ʟ����-��N� �(9ߖp�0S��vH����5�z�`e&������_j��E]��s�<���/�Ѽ���o�<9!I;���k�n�$��	~��J�5�os����'��Yz����O(p����J)�BN��+����iy��4�O��x��OcO�r�lU��'��3)��f��q,O+_z��������Df�{��ŋ���s����\�k����]&gr� ���u�8\y�I��۝�/�
���lw-31��c^���Y�l�kg��L�D5p}@*����'�C�>*�;��;���n���x$z�d�\��ރ�F����迟�p!�w���n3��N�jN�-��q;��--�X������
O@5�O�;�-�T����_�� '��?�ݳ�Z/Dd󪫫���������uV�Aa�S����[��k8�x�F_����B�}���
w��P$�ܾO�La�����KYpt_!v��`J�2V}���S`�Ì9�|�n�dkk����:wGf�ckѫr������r�>��+De�r���yr���ι���oPmz��g��Rl?������(F&8�Rן<y���]�L�P�?����)��%<�n|{>����.V#�u)3��������wc���*���0[w��H\��r�v�7�P⎟�u�x龳�qϣ��3���ll�f�F����������P3���n<<�{�>��j�৷�{��F���\q�o[�ך���0�xD�s_F���dV[�py��p�YeIx~��}L.{�c�+@�
��{�(-�]�������_�گ����U!8�=H�6�,*}��G�¤�5��72u�0��E@QY���%��d����C��Y�ɟ�VL��G����u
d�l�ɂz��FNm<���o�wv�Cf}��Q+��`J�L��I���c��
�����Uo�d/�=�i�4�?��m�;�	��$�ہ� J|�}�����5=�&Q��{�>$ܿ�K�����aݢ�~zN��rp؜i����hw��`��W	uz��&�dJ�^�	����9y0w}�,�ujj[��B�� `�U�@Co�����R?}�յޥ!lV��ى�����N@�̎+����f�N�T�k�k ��ԇ��1��^�R���
�z+�ى��Y��~Tbr�n�e�&x[`��j��!ڌ!+:2:Ҳ�>:َ�l6 �)��th^^���/�%�ZVɡ2P��[{��܌��q����FƝ�(B}�˪ߚ�D�����K6N�m�S�,m)<�Kφ޴�c��G�jl�P`����� Ս�zH�'�����\���:��%!7�^�A��5){	G�ͮ:g54�DI�F�i��䮍�,�s����5\�����>4] ��5^%S��̂9�k�\�/�~~��R\PbmTI4FA'm�`-t��3���˛��V�_��Y�_v��*��d?On��b
p�����f�ڙ,�yъߏ��u΋�0~ZIួ�_��"�W��ɧ�Ɇ��%�����p�&��p)�N�k�\T� ��L�Y�O�h�k�0����`����:��:����$���jݳ1�N�X��~���Ώ��q���S���hu��)�)j�hE(�XF\xc�g��d����I���TUB�o^�d֎��γ���&�4��tB�����q��=�4�D���q��;&�AfL���]a�&���׌�ǥ�����c�y��b��/������'�>Ѥ��kA��T.��a��m���mk�D��޲�#7���6d"�=Y�����I��|H��)�U?��\]���@T~�诞�2l��	>	�7Hє7�>��<
��R2�ܵ{�>���#4��~�`<��eq��+ O�U�����z.�����K�f^5�8�#���0U��}�Hř�h����l����X�M�9)�Qm��;�B@X�2�� �(���ut��O�n�X�SVey�I��x�X����'+�޸�1�%��'ՏBtXW\4��B��Y��B�ж��n߿
4m���1<`����{�0�l���:�Rl������=�b-�;[���� 16��Â�.��=���'�25--l����D:z��~ �t�+{�*�R"I�3t�L ���yo�n�"WA��Lrb��Mw%ŵqS�Yk"J8T	�����TH�uqTYzل4|�V��R�ʷ���N��������;�I۳�j ���<�P��Oؤ�6�	4ɏ �`�E2w�9�M�09&�5$�f� �/�x���AcU0=�KֿD7��Y$�T�,��31fZ�z�����G��T��Y�2����ۇ�y.֘;�/%��+���V?������z��cGPt�vɪ�f���E��^Jn�%���(��0��'�R�}#�x���4��+.�Z�i*N�7����̰�� }Ķ~@�t$j8�uu��s��ot��b����j(tP�
�����v���Y(CM%������l�A<���3���I*0����Ke��~|�Ě6;eXFHX�%=��:��0^��u��|�77���:�;�w2y����R~�}�=�J����/��9�Ǆ�&�:�����熁 U�m:3-99z<�z���,��I�}�3�d��Ϳ�l�D�_Α
��>�I��{|V'=�1�cEsI!�����SLv�=�Ӝ[<<ڎvksKdU�:8x�Ib� �t#I.���v���,���F����\�q#'?l�t�F���e�܋Jl��ȑ�`��JG#4�̴�w�����չ(�F��o�d�bɊ�2�PUˏ՞5K�а�N�� ���h�}����;�d�����
c����G*D����C�ڂ�ΚD����.J��:�(�7If��ZeЈ񽖞�`�G���z���݀$/T���k5Y�h�]S.�k��׺S�A��2��BS�����&Zd{|�@mf�p�t�c�7��Β�Za�2Y]|�kG���#��[�����k�Z�BY��G�=�Y�B$����?��rK~�@�g���]�9!:?���><y"I{��{��o*��l(������9����Z��[U5��m��v����)l5��������#�D[�/{guly����T�r�!Ŕ8Ɂedu$d�֥=Uq]���;���'�����(�c �?�
*��Ř��,����`c0���g�h{����6�J7�ZX�,�Y����Z�`j����/�O�J�B	ސn��NlO�����_�G~9vz�TQi޲1�9?���J��:J�c ��Z��Zk��@����=���;8Buz�s���yk�u�=�5�����2���S�5����ǩ�3;ĸ}�>t�b�J�Q�F���.F̊ X���°� (n����{*�M:�5��G=�������}� ��9����(iQ D��"�-;mu�Cgo�RhV�ߓ�(�9�ü�D?���vNn�̱$*)��k��y�n����ٓC���I����_uP��� |c��W���f1�/�~�@�Oy�W=�tg�J�5���)��Ϻ�=9��J�0�-���	��&ܤ!
�7?'�
^������O�.���X����R��1�ɝ�Ԙ�r�p\_��Dׁ�]ļz����}�S4N ��C��3�T����iL<��Kɟ�53��+G�����}��3�A�����n�2~͍_��ؒ�	��ۓU>e�������t2 ��Ƶ-�9YGM�VV�\e��
I�~e�>�2�g��������tKg�f�R��=��w9������^'��_ʌc&�����pL����<p�A򏧕2hF᡾ӳ?hg�=�����P��F�������|�:��<)JT��QT:�Qgu���ֈd�հ'�O����9N am� ;]�����y]��l��&i�t��px�t���a����
5E����OW��q9�H
<�k��5+h��>�{4�o/��Q�2rR���H-��2��!�;S�
~��f��d�7���ﲲ�j�n�g�
�~�V��+@k�A�駲uX<��gB���c��y�¸ǻ�y��C˴����Đ<0w.��Z8E[o{����[eC����	�<FX��"��3�?��H���_t��/����5 ��ޢ_[V��7N9m��z��Q@� ˬ����� ]�M�����vT���{�RmD�ZZ���hG�9�b0nyp��&I���x-�$�R��{��;��?����7@M�{ɟ�#�i��"g�2Z���5�f��\�d�\��1�pNR���7��'�s)�$�<�5}���ĸ6M��:Ĳ���Ѭ?K��>�$�o�IZ�\��E.B�jw�~�2�w�A�s^��z>T�8�s�.4�RH�S)�f�s��1Vso�`��]�����Zo��[ u����"�b�Ny�M��xΜt(�����P.���
/���T�&,��T�&&Q�O��(�};��fW���NR8�*��~�U��T5�h�p�$Q:۞&�3��c�݊�\A�<#�\��ҋ�}Sܯu5y�m�~�O���I���X�������m��]fΤRCw\[�I��br޵�z�Rr�����L^�*��׍@���iF���^��A����;��r��E�XO	����)S�+��D�,�����f��=R��A�`Y�u��ʊ�cIa���Y>����V.�XTt�Uu4�@m���)�Άh�*���$���t�a��[ź���I7b�|��am745�\!��0�!1*�f؇M� M�1Ԅ(�e.��"p������̢$�n��t�.)��Ϲ������OZ����� 9����SU--m�,��6�j�2�'�������E6{�<bWR��$TB����3c�!���mf�|^-ࣤ�{�yN�8���P��ռ\��ڛl�4�Ɲ�P��c��#�r����#��t�/�u�X5u�8���_0�9��x�tB�)���$��<My�tzbׁm��z��1\��o��y=�/�7͠Hr�������mr�2��c^x��˄.����ܪ[r�:�jYd��
�=�Kj/\��4�|���/5h��Y#���$�� �aZ	"�S�f����a�kT�����ȣ�W�ːj����&��� �נ�4�v�u�_�O
�q�7^ⱆ
�����ퟝ�j�մo�BCE]qmZb����_��0���t���R��-�n��P��Xz�VE�_3{�Bﰊ���/+�kn���-K;
|D_��X?V����6w]��2d+I�t��9��YG�t0y�U1)�W�Z�LcW�l�+�a*d&=�����$�%�������Ը�C�~�T-�+� j-]�L�e���G�/�9e�~��B{���1��3��,��?U���"��@Uq��>ˉ�����V!��~�#x�\��(bk�Y��W;R�xdU7��7�w�7�����CЈ�a���o�1)�܄̺�h֑4�Ƿ�"��)�v����2U�� q��^�~�Z���8tih��
{g��0�����яJ~�&R�3�&��Y�PZ]�/[+x��i��&i
�U�Z��:N�X2��.^����5���,�T7T����&�Oׂ�´lf:�I�f���N%�8�b�@�}�\ŗ3�]�ת������Y\Uf�1�b�k�A2IU����u��K��@�n�Hڱ��)Y㏎�M_��B��"����z�Y;���;�9J$#��%����7�W���V>5=a�@��뮉I��Q�ba?���[����z�x=��{��
p�R�X�p<�=-`W���+�f��k%�ը��8����`& 7�K|6/�a�u��u&���{h�Q�A�C��O)rV�9{���g�5	�]�B����<������z��I�Kܕg ����|�O4~U���Q��9�����*%5U����Q��JD�}�M�ζ~�E�0YB�2�0�Y�"����U3�_��0wD��.���H<��C�7n����r޼�����]����[���b#;��8~ Ϗ���G	ʧ���x^��l�Y�t
P��vZ0R�I��u0P�3�q�I��+P��Е鳓��;e4�R�|��7�)y�n��)Bmi+�b�p�����M��+��b�hS��(E?�W�@�2H�3�f��69d�x��T�m)quw��=rcW(8f��=	��saw�9��!v�ӕ�>���U#!�p��t��t�\�;�H�A���?� �Oյ�~с������ /:V ���!��	�� �M�� ��/:�K����er�	q�o��<��k����ʕ�m�1-�M�;�0��X��)����c�S�$��NO��c�V����,�8^���;TYc`���?I�l%)QJ86J�id��킧��%�'	/	��ǭ�t�˟9�L�p�F�B_�G��lx\��\�ЬC#��$���m'��vr��g�2�؏Lk�i8�a�3D�;;J���AH���p}�d���ܢ!tx����!F�Sv�/�q	I���8B�Q��K�����1��ܾ3����79HИ�[׿(�IQ�a_Ӡ�(��*��B3e��_	gg$a�@ө��4ŕa76nȏ-֙A(\_�2Fǂ�W��?><�ڎ%|-H���4e`�)���������E(��zw�ʿ �ϣ������t:�X~O�zl����|��K�	y� ��ǎj���}�f�Ȫ��9����Wt��xx�z�>�����>	�c�Й��P�4ZH�D��$S�Ӕ�v�L�+��T� �l�; CHe�26f������jH�(�=X�b��~i	I�A5�g}^*��~��i2�De+���Z�:#�g�Z�v| ��w�*���mm�>��]U��
F�D��ȩFG�c�r.���L�v�H�Y��Ҵ�n�$A˅qy"o�5o$k���K�B�m��<}l7��+.����O1�Y����\W���d�ڕH9N?m����]Ԣ��o��� � 6���E�¢��S����9$��=+Fɟ�G����;?���ݱ�OZ@�ˤ��5E�����B����]+v�r��;s���=�37��!\zj�q�!V��Z���� QAxw�{�fv��k�<h�C*hXh_����~��ס'�w�J��ì�Wd[�?�� 1=(�7�g[dϢ�6�p�j�|���ܵM�#��抭�f��e��JKt�,�j������ ㎉�R������PݐFu<(	%����҉��!!���`^��^+_b��/ժ!c���Q8�٭�Ns��P`����X����?��HR�+~��(�����s���ruU�`F�q���of�D訰�hJ�i��'iә� vzVA�돾�e�ȡ[i��n.Ls�GZ�_�u.�eQ�}H�Y������#����~�bͦ{B�!$v���u���<���m��kSe����{hv{����M6'4&F
��_�]�bg.}(AR�����2V�g�Ũ��ۨ���T����4yQ�=��yE~&�[OOl���'._����'輒U���G�k�bI�	����ֿ]�7�Q�F�D��8_�+~hS��>j�n__�_B�x*���X��{��|��
W�G+բ1��䕭$pQ>=,漨m
0���6_e%cbsP�t�ix��	���Z�c.dޢVk�p�t;�����(�#*��Bw�f��+I��8� "-���L?J�O%n1;���O.e�㭓E�}kr3�	Ð养Z�E�]۵�E��!��u�Yl���*/pvd�|�����Uҡà���*S<�Be�Xۓ�@�+�zz\��?�6W�(NB������|�f~Dgd�6��9�-�Ф֬���2�b�;��tĹEl��O,���NI�8ZLH@��w��f�H�4��j(f	(pY,����
��e��b�U���>5��?
�a���o�jYK8:ݕa?�l����l;q���z��G<
8�<�JH����,��!�z��&��nvV/rX��r�i�(�.n��N��RT�^N^J7Q� q�����X����y�c��v�,�T�^rN�F3�J��j!��9(��Kk�k����,,(�G����׫��	��.Z��D���(pPp�(yܛ����h��:5v�;%����\�[J�Y�z��͞��F��>���K�e�+b[z�U��L�������[ぞ[+�78�	Xg
%��p޷i8O��UX'���_
$�+����ιbpS�e@�-v�y�Hq�>���tK/ը�-M�Rl)_��w�D��G���3���� �*DC�dX�i�5�}
�ߑ��ӻv���@�������d"I���x��p,-e+�}�%7�%��t���@�M��3B:����/�2��&[�M�����ݥ�k��H��<��b`��?�3����4ڝ�S�6��/���[�w�2Sr��������i�������oƋ���l����~�M�S�Qɗ�.��$���n�*����M �c��ڳj�2��R*�)3�~�+������yQ�_�з���H`�	���C���_pS�znSƘ����ף Ni��~ee�)>��5�����Lp7~�\S݅ϑ��	�c==2�(4�  ��e!q�UK]����BX��C���#�2q�τ6�1��ץ�y������eFr'��eĔQ.#�d�LtR:�!�t��jj���֯�F�ʻ�����&T�v�K�-A��C�Ƽ@]��V�-u����`3�c�އ}W�J���C|�3e`2��Tw��T�O�����-�>��,򔌝Q�IT���.�[�Y�^�4�=��@$��ɼsk�EV%LɎ�4f4E#�/"�;�왻��T��,���L���>h�H��";�"ՓX�-B�d5��Bůl{�SR���^��h�� |\�?�u�Dȶ�L<Լ��
�%6#�h��he�*��0�VA�DMK�Rh��?1�I~�c�d��a+� ����3�C���m���5]ro�ی����F6�ہ�7��J*7��մ�A�y+��Kd�;�UV��:[���Cv����[-���l��6Y���q@kq�;.�ٿm~�C��V2�TL{&�(�5�i_�CH�Q�`�znx����o}}���'�� ����R������q���Ld������:��r�Q0��L�(�á�#Z�T8�Ax��Z�fߴ���
�d��]��� ����~.>]A����-��7əx�?��8^K�C�	�^d?����ٓ�1Ɵ�>On��2]Wa�t7�v��XC7�%����m�p�Y������K
��B+[S�Xhp^T��v==j	,G5��K���Ȼ�7���)K��� <����;i��R�f��׃`�׵����BipK5���J��"�UW�xee�
�K��L��J�m��'7^C.��V6�������rAzo՗���3W�[����kP�p�-� �/ϧ���|�uE�!M\7���x��8��y?C�G�����7�"W�֢(R�@[�����s�Tt��O�3�o-�v�.����?���c��W��ixz	�j������ŖD�0�V��n���R���<��G��O+�8�>��?J�F�a}ZV���b3Y�g�e�uA��������.��@��X�_0x�������8�tZu���L`;o�f[���_�Z������7�s��lf�m�s
��u�ض�"�"�DF؊���z�kK������dy��0E��(������3NE���F-\�����!��@�K�u�C�k5�%cL8I�w��W[��:}��֕�]�>_�����&��o5S�j��\ƞ��}���*L�X�,���&����W�FFg/�≛��+ywH�v��)����syĖ}����x(�1`��c���m&
�E��5�<�6xgL�����8�'�2�7��kC�C��:�R�u�_C0�{$=��Y�3��T�`�9P��ĀGd���h�'�a�D(3J�.g���q�^rn�}l:��Аʽ[���%Z�#%*�!�~Ҋd_��b�?xT�y�-|���N��J����+e����f�c�#�(�tP>:�_+u�~U� �ԫJ+z7���<r�:�1��v<���1m�.x���'�	z�{@�������)q�ʘq�B<��M��J�H1��O9�"�i�=���^�L`��9��������_�	F�>'?����L�W�KЯR��T�w�ק3�KL����=��ոI���q7D/�߻�~�Oi*p7L{jJ��0�pTU�OMk��`�p�_��������C��H��@V���rm�08s���!��WP��-%HR\A_����h#�6��Y�UR�����#�+e���C_����bu��@��c��[(K���GШ��M-,w��7���G��z�o�N���N��(x�:�}$@�,�%��B��
�V��0n��uBG�#h����\��݈�����zV�z�Ks-�<�QGEr���Y����_�b����(����{�Z	���G�@�263�22]�1�R������d�Q����732N8����yq����E�<Y��SY�B9]Q�6�ua�(�!d+�n��c�W���~jr&8�T�y\���E5o6��0��D��nd��4�5���'@�D���Jp �|[��C媟΢4�8��fYV�H�z� ����X�~�Y���!���G�mO��Sx�U:Da���3�s^���U�a��i�qq�Τ��r��jL�Ī�$܎hT�v�J�g�pJ��J�f�ػ���I�АL�oϻ.h�d�p�r�	��5�j�u�Q��1���E�&���\��N��$W�[�E+���g�n�`�W\؟.X���c�Z7=������^��M�uJd�Bb��{��G[R�9Uڌ�a�����g�����S[b9V�=�$��#Ѧ���CѸۋ�w����T����_��gD80 �_NNm���VH]��q��u�E�޿�#�D����q�P"F���P�[���
ݶ���L����)Ӝ���7�n�J�@��Ѕhb+��wǒ�����A�0/���#��?��:q!�q��u9��o��yH���Z*z���'[arڎޢ���UA�s���hiI,3���/Nr�&-���V!�oM�տeR�ra������fz]���~��B�QJL���Lph��=9�P*���T���އ �ߦ���&��u��Xb#�0u@XلQn=@��kCUV�9��S��y)[������G��iS�6�9��`�a�َF�ov�g�����X��Δht /�i����W|{���ѓ��U��O�`�t�Q�@<|F!j��ڶ>�@Ql����I��O6���yN�
��V,F����b7-�6�Urlڡ��Ș�bl=����2���)�0�)�f`���B�?��)��A��Y�bܯ�W���ܜ�����/�E]�׹�Wu�Tʓl�{yr�.x�����_S�d9�q�	@������!U�lo�rriZ�d���N\��o��j�A
��Ӷ�+y�}���f��.�𤕦6��P���4mA���J���8�o15׷ߘQ{����g��+B����f�-D���TuU��J(��~G�cͪZ��/�Ñ��*�w�

ȷӽ�3#{݇��El) �ԩ��P�I��6�U8�Y��]�Ԭ��u�7O#&F��Κn��x��T��a��Lپ�
j�r3-$1�e`�O3F*\��xk��|1s�j�P����)����W�9k�U��n��)^P!��;�w5w�{�8����ܔ_��=�t�pkm�?��ub�O��^�WSYv���׺�_��l�,Y�ȩ�pK%�U��@���-�PXQޤg��Kv��v&B��b"��Db����ֿ3����ן��X+v]���R��uo����������TQѤ�o�I�Y���O���"z���\��bF�I��DǏ��B�ژ����"-�}�|rj�����uX��]�Ol�o�ҁ&(���\wj19'��M�~�ൗ����{s��'qW���Z4b8|�<J�9<���X ��E0��3>�'D�t�If=���(_��D˵�>*���$�����+)X�Dɓ>N��goN����%�M�t����Ì�i�������`#��pYb��;���D�n!sdij;V�����_u����Ct��7��2��F䳦�4z��K������Є��gXTW�><�L,hb C�ĂR�EQDA@�h 齏�"
QF@� �m�H Aa�(�0 ��9�P�������z�"ל}vY�^���>� �n"���'�U@�ʾZ:v�%?��y��RP��O�WP��֎8`8<����5/�Η�㖜��'�_�a:ߕ��x4��"ںOf����{t�ݬ���o8�_=%�m��a���{�R)�ڑ�F���g�:T��(���b&������M��~]/��HO)? �-eB�C�W_���*������9t��S`���s23q=#�r��������E����M�:�W���d�<_�5��Dj�n[
�����X{&���c{�������%��,�oη�ǁ��Q�&�������;I���I�\H�w���|-@J�I�^�e~�Ț���F�5_}mi-6�'�o5Rג9��ۈ��Gm<�J�����d��x���,�Ǔ�!���ڗ{L7�ن��ʸ����?Z���&�����?���촡-_�<K�(_D��DSO�.��#,�:��]�'X�]����r%��ȣf���88�v��B����qX��PVN9��&������쩆I�0�}R���>���ށ���U˾E��X��E�5lv����������M%��eiE�ͫ�qgG�߁���cv��2�އ_5d�tD	l����ui���g�Ԝ�-E���j�W�*K���`�����.���S�/L[J�XK�d��o��� �6k���b��_��}5����� O��{��ek�d0�mW������=�'^�l��A��F��eo�5Aphg�Xm�0�'*�!]˞[�R�bd�>�Y�-̊z�l@��`�����}���>��,�_ԏ����gfLp�>�%�ī,�̙z�j,�ZA�/n�z 'Q�<��_c��eJl�hRIե���)�0_~x���|���=tl��ޗ�G��� ���]�7EZa��N����}�-y��:`��:[}K�} M�@�N�"��	�f~žڠ�;P���6}�}�4���/����ν�Ik�*n�+q�����=�l��� ']��_\=Gݽ%��/ᨹ8��F��kL�E1��d��:(.�w��%�l�M�� �����]Ăj��d1��fy��l�p�K��2.:�������U�����_�����w� p0o�֧��(Q� Ȧ	�����ꖼت���b��~����N$b8�nT��$�B`����y���h{�I��]��?�� �����A����3Պ�pG}�:�p���GŃ.Hm�8�� 4�F��+	w�VD������oF��׌!�.4H��3��{�|i/�S�j!V��)�I'�5P8fʔ�a�t���n�d����~.��b�X(��_۞����KY�)�P.��{�h4?�^���d��
�N���ehz%�pt?�|�'�EA�;Tc���M>��Y1���"�/�&&ZР�gao���ԋ�Hi��EL�?���DYc�;�f'4�
@ɋe�ɺ}�)�H������5�t�������������g���b���;�<� WՃ���noP<A@i�'��pbq"�jwN����"�[��ͳ�a��%���������]���/׌�����J8�p����K��F�����G9��v~^%�R���+�*;��W��N�f\��,�n�!ע* �_S8z�'��y���`=p(�b���mY����:q�*�/�����:�">}A��˷ѧ^�u��MU٧��4���?�M�iz�K<�~:��]�?E�l�,�HE�.�3�����2UZ�;�}z�X�����Gf7�K�jX����ʲk��	�3ypFx�|-������D\r[Oe���vԄC�L�u{�Ꮏ<:����^I���{(�O�m��9�yth�O>6�	j�~��Y��np�}�9p�0M|^��X.����X��	��?��(�����`4E턬���.�+O�{ ��V�VkBU�Nm��k���3��gW$h�ݶٍ�耤k#�� ��ϛE��޹����g�oVs�����065�0�9Xv#��O��	k�}��9 5W�Y�M�����.[��w���h�\r)�p]F��O�M^ �tw�A"���v�×�0#�P��D�n�m`M� Iz���T���0h�����Ur�HQp6��7�\wo�<�TB#�O��q��U6�����,��znE�_([�G�L�;����ǯ��N����paW]�G��	$ɜ"��%�;��g3~ʓ���K���eb{�p�숄��yW������(H��N�����p���D��ǧ�׽%��_���p�ǃ���|V�P�~��k6�/ݓ����?�ޖosd�5��'zڏSv�	]�s���v�����*�P��ۈw�P/����vן�_�zۉ%�`"Ur��h���x��J�݅I�K�vd��qw6	%�H��B�n���E��˚���;TE@�S�D��M{t<��I�&�V�����F��
����u�����#�J�����A�a
�	���6��N���c���k��k^�X��m#¹kǳ�XڂMBW��{_��_C>Q~/���K�g-K���� ��� �&�r	�G��������fzP)K��;D���A��a�9ɪH�q��|F����O��r��3�,a��3�"i<ǵdP�ZN���Hwp��(+_���=�����ˑ�7�oSqr���dm�+X�T�v����� �+�={5@"0?�+U��ܕ�,~�qy�
�,y����>�0�܂ů ��'�AcQ$]��ߢ>?)e��ζ���uo��,���kk@�� �Zܾ�����$R�B���/Yso��;��D�BN{������2Q4g�/������~Y<B��kO����GQ������ϧ�g߰:��?ڊN���q���ώ5��;��9�+m��yK������L�ܼ���n�r����R�D{������C'/�n�X�;����;����;����;����;����;��B�9�6�R+��л\���^���R�pE��͉K�..����쩝�L-|A�U�v�ԓ�z�E�b�'�%v��7���^�˭���{���{5�ސ�CGVZ��7l������]�#���gҶI$\{�LHw#ZY�c��YI�Q!���5x�H*��n�L����ZH������˓�2�F����H�݉yVf�n\���Cs��"+��u�_c31����1��59g��_К�o[ۚ�E��_K�NL9�ipTCz;6���s�؊U����չ�9�>7��\;�ҳ��h��Qd����T��엀�t*�0�X�Ŝ��>H��A��-g�t��-��5#��5U��ji��ġ}����ڶ��~700�Ԩ=ňgcx)����4�>�0�9����1g�,�,��Ф��ϭE�@eW��n�ų́�w�	��~^�۝�~�`O/�R��k���w�㛨ў:h�����ō���bK������:m�(�AJ��F���Z'�/���G|=N�̍���^&؍��/=7��Ԍ��^�D�@��r3�h�|��G��|�>��a/7�� \5������2�ǱnV,i�	[���p�# �m2�4�B��o!�����	��k��ԟs����;rK�ml����er�#2c%�R���̹�x����&*c�G���a�Ka(ֺ+1����u�-�D���^��v�z�ў�6[�٩��Z�}2�VIav��E�;̍�A���I��w�Qsʼ:��b��.�� �^ݵ�3e��p�թD��;i7n�X�pw�d�o$�NZ�9c�!+pv�>6
�Cvp韮�������y	�I�#��H&����VWt2_:��1����F��3�a$�Y�Q7�C��2��2!v�LW|� ��t��v�;ג���l6k�R`Ppg&d���φ[�:��������S;�xǟ���j��[v���¹�Bn�V�Z�l�dH�GG�9�82��ue�w*C�2O��p�3��qj;����qP�ZN�O3{zR����-��+�z���n�[�F_e�AO'��|.E��M�!n�K�M:Ag9S���F�?am�1�rN�α�8hNJ�_|�]bE��{�n$�������#}ֿ<�=�>�(�����ư�W� ��eN�Bz�F[�#���t{@�����,.sl�+Q�[5|#`���Vy�"�-���=���������ߧ"�=:5� ZX�$"���9�'�{۾���4J����nΗ?~�reB���pe#��0 8(�}��a��֩�وY����~��'�2ݹ�ΰ���7����C���|�餬f�抿0o��&�ٙk���[=��\� �u`7X����k���_�y'�>N�3�v�x�XH�I�����e����GK�ʿy@/uo�����pj�������'�_)7~ҋ��M*�՞{�-ӱ���������ý�䴁�T��G����(�z�c}����LR�@\�j��TK��LS���/p����������-�:~�w�����I�y�h�A�N,q6]�E�V�]����xt�ˀ��m"�/0]�T���70��5��&]��Y�
�|��&N�.9��Ck�mk�����dT�⦾Zց��Dh�E�ȵ�6�RZB*�+�?:W�vs�q�a<Un<�����0;�/q72��κS�Y��t{��}k!�V�/�k�w�St��$f��6�<> �pE�3�3���h�����Ў����3���Cu�[�����F��7�Gb�{ҀF1O�tmT2RʉM���Y�:�����]����뻯�A-X��?-l�w�[�ͻ"T�$D�+��.^���� ���T�����
����3�`�a\Xf9�=�k���و�^��@�*�Aѿ�	?l4D�_��/A��Al�{��!���ީ������n��Og粙�44B��	�@�3n4���jh�$y�������bi�:vƝZ/f�yw#��{��*?#���PAN�ӟd���KH�2�~5��ݯ��OJB�� C@+m��+�3S_��C�j�)��T���{��9T�=l�s��zK�P��Y�kՋ�����c^`�)��W�����b�]5Yr�C�:1%�6,�Ӗ~*���DC��
D�Y�Hj�o�_��xd���!ڿZW���	�G~s��'��a��I��NP9�'�h{�q:�h09ikg!�Vm@�=_��R���ݛE1�$y�&L�nu�3�=�og3.��A7������}v��kx�	��RL���E�I陏�i�0�X O�� Yr¯��1�¹�%��1�P��.|�}f�)����vZ�~�|�Z����ִ�*v;O�6h�vw�dP��5
���t%:�|ZC_�����80����Z<Y�A��e�zB?x�iwGX�7 B�yS�M�{ib�5�7X�@��}PS�K��U}?��
sd��4-���N������Uv��̼߂\h���A����I爙��N�)���ߓ��+0s>O^�M<��"��9���0�;W���#��фi��9���|�B��"���hL>�2`�E� ��S�A#�ؖ-��J������l�U{�#q
u���ǟ;e�x��A�l֠~9l{=�Um�Q��?a����e�]�͙�S�J��NF��D�O��z.�n(��:X���|�Y�M���>Y>�;f&��Xg�+�K"����O{d�ٱ_C����9�0G�m�H�����0ˮc�'m\K"��H���Z��f�/���j-u��ؠX���F:*o���3�
|J
�*�O5~�H��r
	�=�?Q�[���9$H�Bb�هC&��Tv��Ǳ���T���ֹO��c
�4s����/�fm9��з�F ��k"Ǣh�N��(4N�.�㏯�� ٻ�Dd�)��'�Q^�>^�ItJ}�P�;�^:d����.���m�ԯ��n�+Y�4 �#k�}[a�%Gl�Q�v�q�£�oY�REhc��=�q!r�C�|��[�`��Q�.����q�6Ŏ����o�q�-�O�q�)�3�H(r6���Ab<.�A�_&��z��˅���t���&�jBk�ܴҌ�?/_�v3�1���Wo�tѮh�<Y�zKt[��츽�F�3G�T~�_r��2�F�!)W��Ls�������!eR��c��n���p�:.Fa�S�=�/�K�F� T��#_ـ儼��w3�:)����3�j��L����)	}��"4�m1�:<9ܨ��ѓ)�N����Frz-4�F����J���X���E�}oh92{�N�1(����T\}|�6���K,αj��m����E��FUJ]�hP�A�t�k��{|�\�GP>c]�6���J�F�R��q�@n������c�}�{S�Y��pr���0#@ [Ef�][Ψ���G2ػM-L.�~�S1�u���]^�q���hx���p�nޮ[?�ڰ"�]Z���"\e�Yy;�f��<m�Zv+.uB6<���:6��+cl��Wy�xg�JYde��}�I���x#1���O������#����rb�We��.�=�/�<����U������m ��+�+�\M�@��o'���zųo��Z��19v)�P4��N,{�P~��X�r���c��e��ϫ����c�B^��2�p�I_/����©M��Έw7���ƙ�柜9�w�t�jA�L�o�O�3rm9�M1�-�\��NO&�j��X��oOx�L�o:���e0��U�J��� ��c�����}����{��QVME׮��Z����j~��k�\P7��FUM>�U=���6�H9Bp2kcu�*'����6��ߪ'���|!���av��v`�3��zˉE�P���5���i�Roْ=�	�&��A������#��ڜ_\��a� �j���cg��	%��x&n'ì�'&�O]`b��Sī�]�(
�(6N�c���?c�ާ#�9f�~��k<c�b���2~�b%�����a x���oS�bsŻ�:�!�z7Qǧe�{S]S�u�\a$4�Ӫ䔑fw��=cO�ZU����E����6|���
ob,��Jy�*{1-��}\�ݗ���B0Ҫ|�K��u���/��N�G&�;F���m�/uϫ��� �p���5�;�{8L�,���N�*T5ɢ��C��VE�j
?�������p��t��ޯ��_s3@�a0gR�79s��q0���v��V?��ԏ_@�$U�w����X8��3+����}������$o�V����AN������}Op���j)�g��B��������A]Ǽ�;������)��p�xu��H�~���/�H�:W��N({���(���ۛ��N��Cۻ�N��o}�e1�	D�"}6�(hv�ޯ� \����&�?ͫޜW�ܦxE��N����Y~HF��s�֯���;a�+7��\��Y :C��+rW������I'[�����i#��k�g�E`�QM��
q&:�
4�-a���\%a��i+t"����u�	i��J�h�$l�q�y;ӮwZ�?ڱXе���h�,�U*�� k������0?h�%U��I�|!Q��RT�����3	2��T��ɌšMá-�o\��+z`�'���b�Z��X�0�a�O�ݨ�<mzc��Gne�;c�dF����%��
�,�ыQc緙��5��ˎ����SS�bw�5_���R���7w�)1������,^j|�撡4�i��kۊ�9��1x\�o3O �n�i]Y���	��</��99��ƺ�gbL��(ur&0'�?��#;�9�k7�Qp �A<�x�\��=`R��>���beE]����[�2��)1�>r���.��_�W�ɕJ�| =����ޏG��j�f&d᚞�`���CC�T������8�#��t�V2��T�xv�wt�xX�q�KUE'8`��ܛj����!G�i���&?a���{��i},fm�N����F3(�و�]D�:�Zd�>��{Ã�;�	+rf�_nv7��F�*Z8��Z?S�@GI\��xȃ���`��R�&U��������6�8���O9�����5��%!W'���9 "�����t�	��|*���@W1�ZX�f���en\	W!�����Sl>N��s �t[�����M��T޻;��/a�\O��Z.OȞD<��9��0��U�<9�XR8;h���cI���E2�do	�h���D�� �n3us�ޓN�Q�F��)�I��U�"�����a#�Q5<��
L���I̡�����&a	��2��#���@����p��dt�b��w:Gz���8oº=H�M:ꉸ=�+� Q��!1�5�C��n��\O�0��#��v
��Q��+B���]���4JOy����==O�'U�e �\`b�[Mǻ�O'QK���3���P ^=1�JcxL�ĊQp�?Gd�m�wy��nl<��,1U���Hi���&��eW�m@��<e�l��X�j+38�[zSAB^@(�f�z<�]���L-��\y�{���C����M�����޶�gW�Y�$t��]�J�u��o�C5pvƵ3	����!��YeGu~��
�jά�C�*[�;��@��n��8��*L�fv6�(�st�7��{�R�?\���BܖԜ�f�ޛ�:�.��]Y��5��I�3gRZ~��t��������R�k	�j�8n\��E�نǜkl9�<�8hS����|Y�$%5/p~�X=-�d�M���OjT<  ;�;�Ie���	{�um^� K�x��/2�ᕹ�Xc��ԣ�rbc�q�`�ź�K�*O�M��EI׌�%ݻ����C�bT�	���B�vQEHr�Z�(��J��W�Ai����JE�%r���Y�Q?���!�&�UX#�1 �GWd�ťJ�߫P�����<���v��s�\H�vr�N��Tz$�j�&�7���_l�jdÕz��$& ����ح��q���N�o4U�s�qa�Dx�J<v ������@qo��d��NpN*�}�@��ݨ��s� � �!�D<��f�3L&�0/�U��f+Ф2��*�Վ�P����P�������%)S��ݳ2�N��*��XdJӃ��4Ω��z|�%ȯ.�y�΄[�,�#FJ����v)ԗq��M��*���K���B�?r�b��aE�:��ϼ�4-�Ï��l��6��U�A�.*��4�;tŕ�k\��feKd	��?�R����u���w��L	솨��I�������*��:�� �0M��ÿ/hN�����P��D�B���1՝��x/ɪ~뎃�K�%��8Z�u�X1�&�4�D
�X�Ĺ�S��E�04ST�đi
���� �u!��IS���=)rB���2$p[�758�[�mT��1P�����fQ7�O�C����z0����;�ô��?�H����Z�cĽ �j!�(��8��jTUX3��qj�/mHID��Ӿ�?Y� 8K1��0��d�;� ��a�������;����{�^Y�܆�K����Iԓ;F0�w\mFRj��M����������{�Ԍت!�������
{!/<��,���Ow�}ε�����-�9�5�C�
�>�LK����:��퟼��'U�`y�n�HJu�9�l�nX���zѻ�[qOR��2{ȓhIz�hb�O{�#�{�*{�H��ڍ�l��i���F �S����QHX���l4��D�"b;��3���ح�>-�f��{p��ղ�Qgs#��	ĺّ@�|��[��s���P�h���ȡ8�����P<'Qmv@�+��2O�I�wJ�ЇK� }n�����Ӌb�Dj_ݰ|��x@)�^���j�h]���%$��?�L� �7@�g�����l��;������sM�$&�D������������.�<�N�b�K9�D@d��0��Q�Вs�Q0�Ks����t��t��HمF�
P���Cn=_Hf7������=��@u��)̻	��T�E����:�kR��{���{C�#��H����J�:1��f�������T��b�Ԝ:E� eD0��~�U�4�.v����_����x\0x��HA�x���g���Lħ�b�H���Hl�B�������{x`M�Ԣ]E�Q�X��&T�>X 	�?׵d�+��O�b��5Z`�.=�mW4i�Sh��%y/�_UZ�~4)?�~����")��c���1�`|CD%oS]S��W���n8Í+i����N����-��J�����k4VP��M�H���E��`�z#6l�],�ݔ�ک_�����Ǹ��7����f3 �.+qvY,�ǵ��
�b���Ķ���K���P���b'��j2�@-ľV��-���AF�:l�U#b���+O���z�j=r\5�a�c�|U���kP�ͧ9�O1!B�.RHw��Y�T���r��.($Vp�t`R�wp�l�'"��6�\r��]�/�4e��3�$;NW��8�k��E�hH��嫆,�*��X���bJ�)T���7�������3C�Č;>դ�a�#>-�~����/�������L�@r�LS�Ѥ3Z���-!E|�Wz]�g^��A�ɭ�k�ѓr|1XG��@����rE��L4���n�bQ�;�Da8�H�Dq`d�,?t#D�2�q���Gy˅��P�B"SU#��ъ-��B�
�'b�vK<����A�~'�Y�x���bLM�"�p���4�/0�����*]�^��M��:��WI��Y�����9�|�7n���v����PlZ�	�E�)�����J�خh�!�.����u��@�Ƨ.BU!�&߃�g�=�؀#�����h��뎪��>���*�L����*g#��w�[~G�!�q _�O�{���y��!�#���(��]t��0�Jޱ8����Dy4�� 9�u v�W�$����/�&�w��k���,���"Ƞ��P'~<��	�9X��H�}ha��yɱX��73:�����x=b� �mF�?�y}��F�
@-��#�_IoC������l��`c�����GAZ���[�J�69<�ħ�����	bM/����=�&�pT��(�ina��=L3ڌtU��nr���XЄ8`�[TCSD�x�i��C���zİR� �*��s�l?��EzH`��4v!�=^����|�-�(8��oi�[�>q9�13��ճ�*ԙ��fe�3���!�� ml�&�ˍ��V�Ux+%%�8r@r	�K.�/���v0D;c?Ym�?��b�O��]�-�)��P�T����=��u%��h<���\k���㊍N�̃n�<��M�r��O�:&s;}�g'�_�ܧ��*�2�
�7���'�!�A��m�/fԫ���$e9���X���}1w%�I���1�О���Ze1�ʉw5��?�\D�,��!���.V���W�x��'���m�=���8��ꨶpi$ztQy�2�b�u�j���	�������n H@���Ć�T����?�A&ʙ������YC���Ƌ��W�[�7Χ��Id�i��H��'����
�Jv�_�+�:_т��s�N�W߄���2���箻?ps;�f��˞�_?�iX�{]���
V_�> ���"�]1RBX��|+��h_���Q좦#�eT���#3�����Wa���{�K��
��Ox�����9M�R�@R�.ު$9�L��ؘ���8��1���RO��1�e{b�`T���DM������-�>B):v������.	��T�~��t����.bR����g:h_���M1����J^����oa=;���7e��U�	�A;I���l����������9�x���mΝOgC�h����/�@��i�t�]T'�3�Yp)�E�ʳ���T��=W��0[ݱ��g߸��W�u6��5�Q�xSG�����W~���s����ݎ��ݼ^[�D����e�L���6�مOo�wk\���հ �H�8PE:M%g���^�V�~��n;�ݬL�*C��n�TNb�wL�~]�ޘ��g.�?�E�D��l��XRD?3E���B+�(3���t�w��y�a�
�[����U�x�g�;����sg-d�����B��W[�
~+^���b��}�I�DYH�p����T�,��f���=�+^̈��ln+�rg���s��S���f�u7�&��PnqX%��\�H�_�	�j�[�u*��i��e����*i,���P�O�7��(r�a����AO���)9�&�'N8t�e�}%z.���HUU#����O���8M���7{�q�.d���?~Ζ�r��ju�wy�E�<�t{��Ā�h���9#�I���]��G�;M2J[����S����)�M������+	e6ӹ7�6�i���T����In���	cnߌ�g����z<K���
v{�y�2��5��~t��!�hF,t��vN���xk���}�� ����A4r��n�ޤ�ӗ�~|o?�w*�H�q=���&�hh&��Pf� f>eD_O#����Ԉ��}����ĉ��w�!������ښ��3Sّz�p�a�q�b�j&~5������-����ə��S��h��%��w��0�����0�
��������I	hD?����,玳�N�-�1>�����S�Nhq��ʏ<�-��77|�9"�AvIi[�Ą��6����"|W��z\ko���W�ig��p`�gN�Ee�JͰnL����[%�I��c���݀��2�v�����^RzN/`C�qF}tq���	1bV�]�ճ�2x�2�<��)8Uʢ��ȼ�l�IXe7��D���Y�b��8��;�V����kR���ӑM��|t��� ��ǹ'�<ث�����5zt�K�E��������;_R�-0�;�iD؉ن�Bu1��8��tiLb12D3�bR��q�dh��Z�-��w����ƺ�:���^1D��eK�J��4�j�i��qـ�B.�����A��Н\+�XJ��}tH����&�ﴜ��D�JM�4�Q�#�A�!�Ik_�������Z�ҟX�k��5#(~��V.�=q6��D�X�aR��7�l<.<s���jeg֗j�H]�a��a��S#e�m�����Giq�{��4�gΛ�|��ȧ�8�5�]6�O�H�aN��ե�F�iF����){<�o����'Z\���8<%��L%ݓ�'��G�)J�(ă�NSN���s�kxs����M��2�_�RǦ>O�̊�3G�JC�5^_������7~^��S|�A�����hj|8kب��N_��i�3x�>^�ӕ�<��W�y�2�a��cՀ>�~;u�ߎ�B11��85w�1%�k���z��-.����q��x�@.�7c�}��P�0�����\t�_J,���g������Φ���~���ZCӭ��3�[�$�f$��ˆm��S�2��
	G��g�he�uk�?�.oz�<e��V��Y�f�}�l����Q�r����Z�9�t�ԥC���:5j~/��Li��7��X14���N�U���8K�l�����a�D��^޶�ja�z����Ϩq�Z'�Q������x�0���,^�{��>W1.O�s�3a�;$z.�L{sB[�O�]����Jn_c��D��F��N�c���dn;�s��i �$�]�D��t�3?IMm�5����'�V���:�C�b��u��޳O:��f6��Zd��C��E�*UD����\e���/ic_��#��������W�w�::n�S86����U=�[�`��M����'nz=��;������Ѭɜ�U[Vt�;+�h8*�W���6C/�O�Y�ki��y�)5z��H:7zK@��~����sgL���)YO�<ҽ�
X�7m3҇x�t5b���g�H�r����x��'&AP��ӎ<����TƁ��%�[��v"xؕSy�uiI=%��/�IQ׭���7U��,]�v�_[&�N[�j����F�&�;��]&���}��T�͋�g�r%�^����mf5g���҅�6������p��(�������2z��_Y�45s�7�iތ7)����`)fܙUV�|v��=j�it��v\�C͏oj}_��v��.���Ok�{L�59k3ئ�ڣof&�x�g��y?�Ꜥ�^��qj��.ѣk%����]u�<�ˣ�݌wО�i��%r���܀���	]<�n��GT�~'�'C�}��௉�Y�NcA��p3���l�^�?�G��Tk��Ӗ����i}u�W_��}ȇ{�K/fS[�^Td�����.��gƤq�i)����6���O�ǔ�jA�v����x`��
�F����w��4�׫�L�Au��Z_�TI�[&��{r;����C
B����i�dٴ����CXu��)f!.;vX�n���u�W�a���T
%�A��0B�mmu��A�|R*L�+�흖g7B�QӔ�'v5	&V$�����ĸ���P|Jې��N�9���47ϭ��B�"82i�:z��q�Ln=1��9>pI�ً��A�ͰS1z������#���Ǜ8�P��>x�X�t��t�Ha�Lh� )���#S\ǈ��2�����^Q"�˞��1߷�޼�����	��}�.�Yn���%�^��d��FI9ھZf�ս?�oݟ��1%�(jk����w�sN��Z~�����HuM�!���X;}BB�Ւw�?LBѹ�xV"q���7�.R_&m]�	�z ��J�HC��f��g_�cB�=}�fH,�Y�;nS���`1Z����
��i��Qk�m������`�X|��c)�8RtM��M�D7����qW�6�ԫ��;����d�ѺO��cv�v*�!X�}�����>m���c|���zeǌ����C�Fx`�@��� �3��Rқ�L���O�T 7�e��@�H���j��,%��O���wN�􄑆�[J��ќ��8_�a�vwS[��r�� P�w��O�n$�G�|P90t8:�y�����׽ 8迪�Ć��!���;?��b�
i)���d�Z_����1�r�T�i�pvӴ���/?�@s�[�'󴴟f@Y��4�G���hJC�N� 8��Qn��jd~����0��gM���!�H�6�ޛ�]w�y��7'�#Q�J㾗~�U+cf�|5`�Dt��nN���0�� ��j������@h	܉>�2��{�ĝO���c�-���k�Pa���� 5w��B���9����ѓxG"����a�~�l����X5�Zp���>�$���'�b�w� �~�5��w�^�72N���r��,�L{g�� �Z��z�%�N;Ih+��M,��5��ZE27�B��͕I�hH/"��9���t}��b��РbJ�y�'�A�ɣ\эJ"em$�'��!+Ox�D�+�x#���m�zQ⸷���i�Lþ���<��~�0��U����P�*q�+M�o���*gAOM<mکA�Fm
�m
GZQ����}���#��=1u/B�x:�L���?��)I��CYA�Z��:�쾮����9.�Ȅ��x��U�iڊ�R	�|�$��:� ���O�6]xo�߸�Ï�|F�SYF}��w&�Į�7�N����XW?�&����-���w�}|�9!:5tLc�˭�4�3:�DY�X�OSs���d�z8�(����@�~Y��HiL2D�j΢%��b��΋�I[$<Ɠ����r f�o���M$����bD���Py�����C�r�x
���ף�� O�~/mJ���E�'����@;����-��jmN�į�B(aH���V�2ӵ�Z �:�a48���c+n���!�d�n���WD�_�E>�-K���S�-�:Ϛ��-�����	��(1��y�S����bP[sZ�}"�Cщ"��wL ��w(�`�0��o�~q�L1~e�z�����i�𴓎"��(n^��%�S'��_�<A����\�Ͻy��?Ag�ヱD�A9�^S�G�:Ju����RPұ=غ/�/L�s�����L��4�CM��� E��ɧ��������K�o���PDhHޠ�'��|��Rb�}�{,8�~s�wG~��g��Vd� �nRp".j�麙�ŷm�L��ks���������o�)_�t�f4Ppx��O�D�=]�f���K�H�1;�b
�y�|@b*����r�Y�w��\��������!)�Qu�PU��Cż��:�K���:k�?a᠂�
Q������m��[�^������oy%^��ﾚ�Šzg�h�_'�����b�-� �y9��,��o�[�͖H����l�·#-A�ߦ7i��9H� KE�hj|��?/�?H�]���x ����{��i�Sa̋��_!����J�R�߄��3�(�/�%�
dI�f��/1h�3���
'�^�b��1���L=��S�C�Z��L�-@]�F�o��݀S��8EmJ��r�nҳ����lZ��B���1y�cXM���A��qn�D6
O�CK���䥶A�]t�;������߇*m�"�lz���ܥ�/)��׋�r
DU�� _|{��?j�7P��+7Cf􀄅�HT�]����4��~�qM�|R���2
�����P�� �-�zu�3�a��х;�y���-z�M����QP}��Eڀ'�������$;G�d�_�X��A�߰V�f���U�Η������2�.P:
*�;�%��I�˨٥i��bZ��X�Vޠz_�r�K��6��1ZY,}�#�H����c��]w�3����	R���/5s���?�Ca���6�b���%^9~^.Jغ���-��K��1*C��r�'��?��d�|O�����G�K)�F�'t�S��ρ#-�ߜ�!{���9��ȇ��(n�)WE9�6d Q��"!�w���ŏ��!�Rɞ�~u��qv�¿�Wr~�^�?n��X�4����Mƙ0�D��Ma��죋���p&5w�Z>^X����.�

P�����Re�j,�;ӘX��`�1\M�l�p�ͥ1ʙ�q��czm��T,]���$z�F�tN�>�η����R�]_���/�1��fw�\xUzTN󕓩4�=��Si�2�>�L�E��  �$j�Z\\d�kpL�S)��5�G��&q��%*Ei*H�<xme��+���vI]����Ћ
��n�D!,���|���X�XX3�vo@s-�׉����s�7������C�D@�H�
[?�G�giP�Y�yq���Przs�������M��:N��2�`�b%p�_�`�1����P����^�.�uH?�����_͍n����Qvs�m����HeJm�<Ԓ���W��y&��*���XH5��x*s�:�v ��u/�� ���BA�f�ț��H>&���"�\�[��6C�4�_:�8�mn���"C�8�V�C鞎�AG����E�dSp�sl$j"�X7p����X�!�u�W4j0���SƋ�C�t�j/pHã/���'P���?~gR/���#(�τKǻY&{���9�C�(7��_W��-NB]f.�X���O�4�ƧF�,�	�#C�	�>���Ρ%5�6ɋ���.�_r��K�6W�6�8*�ӏ�[��c�&��UK�'��y�]H,�� zb��;��b�a}[�ԜG-p�z]��~fڜa7e;�C{q&���s=7�-7�]��ҷ�g\�
ϗ��hR |�0����#��6�A:�Љ��#f��YɊGޝi���>.YB*h�g&�vX���D�
7�3��+�q��)����y'$)�4�{�E����`L�Ʒ���26;����R[��� ��Y��C�ݣ����RB@��v-p��:{*�4���_����ct�K�-q;��Kw�UA�D���ʎ4}�?�� [9)(j�JI�	 !`�.��i4���MJ~
�/-�����e����;`�f}�@|�Jm/{� �]��Y�H?��7��q�  H���־���7�H�R�Q#��.�ɲ���2G�=�z�ͦԽ:�/�@?��\B�~�j[W�Tж�$�3dnKpϦ�RNH2��¥~�TS�q6�>9}g��;9c��浲{u��3�c��l��)�P�s�~>7�J�͜�-O�z����{���\.�&�kw2y�����/��*8�?��>���G��?l���t��G���6�D���N��~H�����<���oKCy�5�9ͶMu9j#&H��6�FU���Q;\���(^�>+�-������i?�B+Ruͧ�I���X�n/�e���\�k9U.�yin{]3��d����D<opl5<-<��/$K���'y
��-��_@|��vU+��-�<,t�v����{��454TO��+��։#�Ɯ ��'���5�C;����(�*�v
	U��_p�/^F�Թqk$��
e����q����/3 eD�9���f���d:vZ��m���;R���}�]^�9դ�^Ȥ�5Ri�r?{�#�jؘgj��X�ˁpT3{5��|z�H��qenZS/�9���$ˁz6M�pL��ܸ���nB�\����N5,q����V�][q�vu%8;{���%d����bi�����^�J����ڋ��~(4Խ�x)�2�J�quLm��v�)Ԉ��`��^>��
�w�;��m�d�t-8S&�~�n�Ƀ5��E�>"? �?���%je�Ԗ��:'�$dHW��Q�N��>�:�O���C_�xb8Y�n,�q/m_Jb4��>1����R��W�n�ժ�N�4���[�p��<_.|���_I1N�zҨ�����-�UW#���Dee;����\�s��`m�B�������yt��qm����6�
YөaW�N8⹌�nj<|�ʧ�M��T�.z���Aw�n٩S��Q����V�G�V0�n��»�����d���T�i{"�;��ߺ�t��b�͌#�i�Ƴ�ۺ̞�H�� Vn洞��R�K&����ǃ���MU
+ٛ�D܃�o� �K"�)�c��4e�<%��p�UUd�Z8b�:�1�%���<c�[#��������G���<c���ItB���E�*�u�����+'\ E��磞�V1���.q0����=x�ў�����og5�yױe����[�:�iI�9�$��)���(�ˍ��~�v�9dB*j��v\S��C�⪇+ﺪj��ƕmn,�$#G�y�� � 4.�m����0�sa�2RvPU�X�k����<�����:G?�p�����<=��<�k�<�87�������ҫ1�@Ч+���v{��ԧJ&�{�y-���[�[�׻^;��%�X��~�s���U������\k(^���O�+)Ó�����J	6�0�EՃ�I]/��o��z�	�4�v��u��~�#Ovq��?�y���j|�S%M�;Ŷ��9uD����1]BjjaV�sB��(y�!G����x�0{��j#�� {�m�O��nt*���B�˼S�5������p���L�WӦ	��"�r6��"4x�����������J=���)��T���Z(2aZP�ٙ�J�Ǟ�bHJY�T�^dO�=��;�w������>��|�����?�Ϲ3w�E����s~��$H?t���b����3p͠[�C|�R�n&����ϗrf����#����֤�Y�'k>�t[	E�i�;k����{o���z̶���LG�zx��3�`3mQP�g���(kFڟPQ��{�=l����E����uLav�����w��=E|�\���0>�V��]��� t�>�i|RQilŸu^��M��� 3��5���H����W�Z$]���#�{:����a�_��.�S�[��'�L��� � �ׅ���t��^7/�P6f��Q����|�Z�	�/-/zn�N�y6�a!���`�%���}N�
��]x0�ňP	���M˛���~����ԭ�bD��|�����/"�#>�[S��7�I7��v��l����l�^�d�?`���J��E��S�Лα#f��y{ 8(��	�_�,�]�B�F�۶B��c��+�ߌ�?����<h���z��
�u��}~�&�nI^���L�٣U���ߚ�����s��RS�I]���{'ނ�K���җ�i�+�A����z��Y�:��C�����	%��w�K��kv����h�0��	T0�K�\ҳ	 ]R���)���ۈ��P82���#\o��Ex�m��2��z��9SajT��_I��m�B��js{��б�[�?�����C@y>?hzlb��g�U8y=]�T�~��<��	���u��B$���\�J��,�gb-�y��0'o�j���O�$�Љ��~�u� X������'՘���|����'�г�b+�XhD�)�ʯ|QZ`�Y�� K딓�6S`���LJ�z4��Lw�8�i�XRC�yQ�Ά�l����K?���c+;#�$��y��A �b��P��0%%����������AI����ATsQR�&A���K�[���
 ��S�EW����l�ተ���:�Az����aM�b�����^Iv�У�t"��&}��X1��o\�Dd׽A~P������QK�xE��G q9�6!�+��V<~����&%�#��S��<�0���a��6�]i �`2��2P.��Y��j{�I%F���Byվ���]���͔8 H��lR@ki�y�y�!󋜚C-��V��t���>�e|VR�yh˹R�x���w#"���<��<�����v��7�$hӍTr>y�_R�t�?hn�iܫ
,�F��5�q�4�V�l�Ƣ.�U&+��Y-AZ�7��F:���6�_��c^1��u*J�x�z���V�<M��
�������!�S����Ψ���/!`\u.,9��`�h_����_�";�K�}D�|��E~XNe�ê&�������T�������a�N�-�P��v_R\N��ܟ���e���
R�r�DHG`&�oJ6u;tTt�=�&��+�Η�@��}μ �g|wV�3��5��x�����*P��¼���2�%)3VC_������+ѹ�AMKa���s���2t��7Yee-��f�և_�bL'~�SB���ڒW~�*�[�`i9�qL����ҍu�b@�;g�j���#��쮈1;(���-lc�8)������\�N�aj0�OJjKYH�\�B_UXL�Á��ϧw��r���N���r�=�(("�u��k(Dm��b�K��N�@m'*m]EY��TUk�\�?^ԕb�?��X�{�R���+�FX�K�Sk 3q]�?D���`��T.l'@Y�dc�q����<4���m]�=]�+�Ʋ��FV	+��\lx��3������l��$~��4�I��@�l����b^N~Ԇ��1,�z�W���1Y�hl�j�Y����E�:�V���y��?��	���-F�y�A�4�<޺3�ﳟ��W	�^5^��;��`�l`�Y�	���?������y��ZE�9c�)-<�f~�c\8]���$|SE$�\�>k��#���PU3����Q�n����������A�S��BcQVh��I~�3^�4��5b|Z�~ �\c! <�e���p���R�������C�O�~�9IM�0_*+��u\���������"�YյH�!u5Ξ6E�|�Fb����"Ҙ��{���%Q7��ձa��VBmL�ɔ��MCT�0U���:�2|m��' ��%1c� ˵+>/���ޛ�eU�1���vv�T8��A^��P:#`���N ^�R�*�$� ��?ő�]���/ރ«��g:�[�u���sm>8 6 �Vt�"��>|
\��&����l���m���� ���U�ٷ��Yl��2��P��J�٥�nE�*��ف���	xRb&�.�@З�/�
qs�cR��H�f��������V��F[f�.m��'�C�1�m}syq����d�*X�y}�n�=v(����ї�	*�+Ũo�,�G���
�U��Q|D>�_�{Q�x�1V�#�Gٰ[R[��]!�����<�o�y���&�y��K��o!tN�=3�W�,�]��G�������|�*�����,]�equ�����WvhK2�8��U������ma���9Kګ��g�m��̍����DWn�J��f���0)��\�S�mR�u�b٢���v��L.�,}�X�`��_T\;�:�`�X���%M@T�Z<^U���5�&~�\���@�F�*{��nK%Fv��7���1EڻO�KP��7QA������4�ڬ��u��>׌�L�BM;c�5��|Y��Ľ���S�F|!�"g���@ꥩP5��3�vn������ro�g��,L�,9�DD��l���>�}�i"��Ce��N���٪�}��VPJ3�A<ѭY���ߩ]�	�����F��l�oG��w�i4���x�*��`�!I�V2��Ï��i&�5�|�g1�t�5]��3v\=�#�c�����@��ύ�E��hV��sޭ̸�g�nWqWūY"3)m�qm}���*�0k[��lB���1��=]i�*)���|)�Fti���Y�����{s����H:�ژ���l���/�3�L�����ըx"�
�?c��V������_��psd�uy$%�׫�W!���)Lm��C�s$%ň��}�q��<z��y�^��(L1zl�r�ӕ�� ���ۏ=%U@�9����m�הּo:��$�Ի�����W��uд�����a�`Dy���,|��8����M��*��cIW�0��.D
��r��"��Ct]n�<ba��cq���8�1m�yܭ7�L<�C��2�d���(�@�ׅ]�In��f7r���V�+v<\�$H'��0�י�[|�_�/�z��78�#���=^�T��ű�aˈ�r���Oa
-\�1��S�=�7Mu�N]$t��M��n�K�]E���̂����C V�o-t-wFg��\ي���I&�c�m���=fl��A�|;���/��ʰx�̈́�+�G(zDZ����Ʈ�!��Kym���G�7��%�"J��lw�����^�,Z(�ME�	���c/]J��I�DX��:p6�p"^}�[��U����a?�����u�[*��.�+��L�/6��ի@q_C���N�`����=J�7�_r�j��j��̎�c�:�������Jj���N���"n���;�����v.F�K���FW|<��K�W���H�}��:���� V�����&����HXGRd��-���m�0_���HXF�)�f�M����kI1�J]��;�w���u��T,ў��n Ԓa*��! ��7��:Y�ԧ>s�-�u Z�+��n�*>nn����v��	 d�%��K�h��ߦ.�l�t��#g�I%���*C�э�f˖��4�y�6��iE�ϡ��w�^	cB��C�V��O�ˋEm�9��� �7��t�>����9�u�����A�Ins}g��������`�С�R�8�&p�҈p��qхhw[?t��io$-�I ��W�JxlB:~�>��oj��~��6� 2T����O}��++�6�����m籟21��U?�Բj a�^ځP�\"�Ah���&�_��*��u�\��f���=�79��b�W�T��֠�S\���_��]h_������b !��8��j�@�Yӷwƺ.qx���;@h�G�Z(X�NcTI�l{\2�@�4t1?��y}��y��@�Dn������N�I[�7�i���h�z���/GPO�cߜÉj��HSI1���,�^�
�ng�E[Q/�ڴ��ϻ]�[����'�Ae!�{������nQ����w��iIc��F6�gj�H%��Hsݐ��ב���> �2 ���!�:�FR�Z��2?����C�Ŗ��� �>�K�G"�G�$�;�����hg��lz�]�d�b�]�6a����c��KK㖋�Αˇ�E�j�[�c�!��߄����Z��ŲZ���FƳ���H�OױE�#F����b����}�_9G;Ń󇾚�Q��ߚ@�IY��mU �2����yhK+�!0�mv*c���e�����A�?���!����Nי-�_2���cCҀ�{w�����+�ed��FI_�B2}ض8�{Bj�)��.OVIB�=W�gO�5�A�L���o�vL��/D��n�c��t2��^Vk�E=I�n��nש(6um�h�/z���>B	2"�@�,Tpr�\c�#��ʰW���$zt*��Qנ�lfatO��7��&���G��gl��|���M����pb�h�Q N2-M^B[��T<��KP���B_?����y,�t@��s����+��	��P�<���j^0��#Bv���_!���ā˂��K�Ϡ{�a�M�Y!g��=�L�ʼ�3_����& �m�}#�6��,&@2��*˘?�����-��2b�Q�HghI � @^V�j���D@���ר�)���_�Z]mD p������ ��sϰ4��µ�����+�s��h�/pr�)zч��1RXɎ�p��KV��^+�"�;���ا0�ǆ�n�p� H��c]r1���i~�T6{�Ģ����☖u�j+#��[H�aç�OH��譢x�\d���Ø�|^����<M����u���s��r�}��~�[ƾ`�E�Cf������k3v�*�z�t�5������J|�#w��b��W�4���>�g�3���w6b���}P�Of�������mOqX]a�^�o	4�`�⤹/J#&���@F��:	Ҧ��Hv]{ꂲ�M�����0�s0�?�ȓ�nX�ex�>�E�j��Ȳ���ai��=���t��/�Q�A.~PY ��i��3�FK����j�a?��r6G�FE�lފ1�����'��n��>�Z�e�LVB��������Fg1\weɶ��RY�6�L=�6��ʖ�D<F��Ff=�  T��Ā�#�@����/z�z���T͏���^�V!g	��̋��d��~�"1�np�x�q2hH���ԩ�_��i�$F*��όD|NWx�<�Ѯ�(�L⃘��F��񣚄��64����r懗�W�
�:	����- ��<2�i��14��[��� ��~^�Mo ���@��O���1�_�|SaO���Q�����n�*HRؤHS��ѕ� �G�[(��]u�E?�컼���:�?z8����.H���הF�ɕ?ڷ%Z�]���d�`�N\&�`�&��ғD�Z�FP��ʵz�����W�t��!/یZJh˯��+cL	�+{-�]9Ni�������!�v�./��
D��T�����a��@h&�ۦ�`j`I��z���%�7f�&z�k�b)���}��| L�H��ň��-�Jl��x�LIf̧��'z*Ǐ�.z�����?1�C�o��>�5�3�4�E|Dq��{�Y�C*��d^����*�F��d�		�%#���\��J�Eñ	G�?R�g=]����%�����ư�L&���!1����spf̷��|�^�m���C���c�^2[F�VF"%{�9#��)'��9#��h���/���PE�vn@��t����_4+�W�sd�)���M���G�	-4�Z��í�;{��l8�щ΀������~ʄcZ�݃\f��c�ܠ�]� �lBtY�^�1���C{�{�2�3�.��j���jYۊ�+=��!�/A;GS*��*��Cdf��he27��yx���2�Z�6���k�G�g�Г��x��Ht:}+u��ؤ�/3��49+�Q��V�ѥ	�� tR1�0?{BF�|~��̮�w/-}_F:�6�����Fڏ�R�=�pD�7�����n��=&X�r��G���B.F�`Y}r��K�v0oy��fgg�FR�;?O��Z,���Z4����e��6��q'��-M�7,�H�?�+�
H����{1Y}�z�o(5�׉��~�XB�Z�j���y��x��2Ԁ��P>Kq]��_ rG���t��xp�_v���d�5t4p���M�[�(+�����]�F?m���6y-����	�R.}�˷����(��6��zKz�� 鮂�<Pu5+�=)�ȱ���X�O�/Ͻ��8؝��67�+�s�`h����ݎ����#�Y�@��3���zt�\Ͽ�3v��_��~��[��%���@U��<%�ީՖ�衡�X���H����	$-+&��1<Z�I1 $��s�m�M"y�L}�����R	7	�_��2���+�yy����	�
8C��h0��b�?� 擲�b(̗Z��
P�YEq�!ꀂ���������G���&������,���XVAb���t�c k���H�5}��c�!�>o��@��Bep���E:��@ɿ����S��>���Q�4 �H�z2蟕�;��V�!�ד߭����B��Ձ�r��ͪ��W�@�|N�y��Xt�#P�y�J��Ϊ����D��\�#4�|t����F_T?Ot��̅�k �ߕ�)���dI���'�V� X_T|���2.@��iڎEר�����a����EK�3 �!ତ4�+�uk�Ľe8���{��֙���#��V0d� d�]�����t${Z��:���^MEU�[�8un���Xs:�Ջ��*.�Ry�"c���}3�����?`Tb�K⟦�!�҅��x's�c�RoH��.jI��,��V����iԭVA�u��n(�=.2k�2�\�:T%<� ����|������q���]�Kn
5���|uR��������!�X�Jg߳��"[�󬚽|���]Z��p#�z�.���ֻ'fe������7~�#I?�*/�0l�$I�s�G*sZ�ж|�/�mz����w�Tۍ��3�@P�*�q���|���f�h�1�_��RCR���d�ze�~��f�̣��y]I9<a�zX�][�gq28�m���FP1��5��>�W\��O����o�߮'ޏ0_Z���e�m�I8=TV�9���|��X��O��=��s�삋'������6vL����w����f�]�Y�P���e�vS�'ob���+4��u7N���uZHɡ]�� ��0XX�Ǡ���,�ʙn5}K�;,��M'|�.ZD7���l>�K��+���45���Ռ�.EU-D��!���ϟ�Ħ������h��u�<km'~��W�g�_b�r(v�uZt��歺��D��!W!Ϲ��*��ے9�W��f���G�q�!��z,�~��~�k�_�o�v�2���*x�^�Un1��\A
<p�Au�O��&�1!��]��!)�̙�s8$1�Z���˗���E!��_A��ӧx:�?,q7R����g�Cٗ�!��5�����{aR�e֢!v ��>'�:窫p\}�6�Y�$�hP���L�/�Q���r�쁬(��i���(�e݀/{[ߧ���6��2-�9�.�@�8��l6t?��TM�.?��|�yb���بݜ�'��:�e+�i���o�O^���(�h�'dP����6?�Yup����l�%�v���<��ݚF�K�}C#����0L��)؊1�ְ��2�t�!��3���n[�Rt��P����x�U���(�-�����F�Žߩ��@�.�DbT�=���R[�(b ����G�g+�� rd�A�6bʿ��#��sd[Y��p����@��^(s�ݰ���';����ӕ7i���Z&]��e����c6�L�!L�7�c.yu|�K�_
�IpO8;H�&w�RR��]u���.i@l|{��^�l�Wb�ǝ �*Jxա�=S�> ��:-�Hd|�A�пX���,���S�n�u��A���uT�"u�(&z(q�?~nz�,��|�`�⠽eXU ����w�,�x�G7������c�`Q8����|���huQ���g��i�8��o��� Ф`�ԋc6[�����&�l>C�����&�\�ͼ<rIg��qK���u���c�=U�]W�θ�������X0.���Wn�t��ݜ��(���z�����c�K��:� �������}��^�q��W�q�$�+ƽ�֨�OkM��i5��F ���g8�޼}�0��9=пZ�Cj���;i��������)-����� �$~�H�)�-tBr+ Y��̟��3��1v�0��i#�Q8���[�7��F���o�V�cA#}�����e�6�.�4E�X�� ?��1�MwD����d�O�]�^[(�����[�+����Zb$�S���q*�˽=j�(A{P۹F�v��Xi�,�c��ҡ c�f�^��ÍP�W8�im$5���2��rԄ��rY�(���A�胚Ex0�=fC�����2��¢�*�@*SD��ǴjE�Z�`��W6pV�N֫�-��~@��,y����i�U��W�4�fg|���E��a7#A�6���3��ǚ�c�u�q(��sh�F ��x����j0���5�9��|�ҵF��o��@z5x7'�� ��߀K7���[8E���S��r�%�cV����UK��s�����/��޼��r{���`��i�s�(�n
OԖןb��-e,��^
Dmp�1��؄r�j��=Ke���r6̨�wXy�%����8�9cQ+M�� a��@�����!����� MB��0�3�n@�� �������\L4���O���	� `�L#j�oO�s������1�X�clP�
�~���j�� v�x�R����oe�{���YQ�{1��-� Ye��N�O�)�F`�O,?�~�����sg�².D� 3���Qmr4p5�!5��dX�Ӥָ�F��N��%b��;��jB�h�;Z_ؽ;J5@���];ʃ�iR�5��@W�X��Z��^��j��W�c�é"j�G��9 ��2Şog�.�J����l���0)�P�r- Q���X���XH櫿?���&��P�V�RV�4fz�>KY[Y�Pbݺ�"�Ŷ��"�|e�8��o��
x2��
~H�4�!3k��ӣ�Ig��c���.̽�-Z
Ar`k����OB��-Ɨ�����c��f�3~�̻���(�墱�k:Q������&
+.:�?���-C�CGD�7�1Q�7]�Ӿ`���m�h�$a���Z*�xr.�d��
�|r�O��̸�tb�������:w�[p~ ��|�	������B�n��R���F��?�,M�حE/���|�h�7��A�e��٭�_�Q�#6�{�+���D�}��l:&�_8M����� ��y�}enڃFY �liU�~q��򩧫O߈;��r������Kο�pC��kL_V���Ő�8�p�3�3a�gZ�g����4����y�:Y�U%�E�7]{�ia�5E�c��y�_Z��D��w�ȳ�@�|�^���Z�M���S^�h�ݥ�|%�����c{E�S�_�[^RC ��(�,h@j8�����5��X�g�' P���qʓ�˞���Q� ��Tw��\�N�%K���~�E�6��c� �.��{������j*�G&ت ج�����d���1S9ț+��9e*�9<�.�,�N�ݥ���+;o��(��e�|r�y�L&v=g�f顆��]�-K(ڂ�*S��SB����}?�1�
`�z���bI��R�!ȑ��8q�HX285�SC;KV8�%`�9���qdl����5���J��+`�M=ʳ��/������=�Fˏ�����%�<	�*2���x���[��b����O*:	�C����m�%�4![�;����-�0Xt��P�iE�4[
H����L�}�{,��~�!n�5(�җ���aO���Г����$�
�!;��U�\��e�N`���Z���'� ���:�,�!�zNw�_��<��>&X�:> �;�4�N��}>��~��Is_���/|t�1��{�<��W��p�*������vtk,t�x���]�c�f�;��y��1O��@�'��-�8���-c����*�oG��4���M
���>FЇ�� �K�h ��a��%���7r,BZ�K}~0 ��z�$0?��q�_ve�94Z��X����+�^�	���3rB��z��;n�V˼���'f�&�&�m�����3K�7�i6�ԝ����������h��,�LY�w��dA���N:Qg?�`2O$�H����M���A��N����0��:���g�P��V-��6��i�u�0�����T.�AǗbHf�{�a&��Џ5��kӋ_z�%: Ё�������}Q違1��˳���d�p&n���(�<3����B����gԯ��՘�Eۣ��O&z�M�4����f�p&c�dcy]�T0Vy��!@i�MF_�Ͱ!�2	*Y���+΃V>�F0����'�5��:Fa����5�7z|v��B0ܩ��7���6�X�=զ���F� `h��o�T�[�(�~m~�L�߳=��;`<�\%E���-@� U�(�O@C��~��S�?�`�B��??6R3��6 �;���$Ւ�߶u>*���W�k���S��ZD�c��:��"*�SUI5��)m���3O ��;��AR��װsz���1 �T���K�C=��9Mb�ƅ���|=�c�;��y�{5�<�~v�/�� ��O������@���n����3� 3�
D�o�}	�0p]@]o}c�1$��Έ	�򠁜gҕ�
���X�j�s�5�H��e�s�Y����`���r1:���m���:��������'p0Oa�ߕw+ ��_���C�#_amZ�6������쵹I��~��اiȶ�
 �\�*o��g�[w�Z�9�,���_XII�B��l�T$���JnLZ��rꡣ8R�d��:�[� ��a���Pf� ձ��_4�$�<`֬:�aC[,cqp?g��p�Ij��}�SC0��Q_����z�� �������>���N�n�/���?���%��W��/��|!VT!VH���½p�s�F W6�����x�/ڋ�����
_��Tg~��,�w�Mx$���3��<��Q�k������8i?$Kʱt^�`�;cM���1� ��P�bS����W�)`�l����1T� W�f]T�1���@�m��x�g�5����U�(T�g z(�/z����X�Z��B=e=ق�D�z����S/�2n�j3��YM �yβn�ڹ�C��t�(z��	ڝ_�mcX~��Ƽ��-�@ka������&���ԇbG�������6��X%i}G�q��D6+I�s��H|�z��H�ʃ
?�_
��	�1� �^�v'wn6Ⱥ�ȯ�����
�� ڳb�AI�Nz�/������?Agx���40�UI�d�z���Q�XzȨL��X�:����=�Ҩ� pe�t���� �{���`����<��4��:�[7�)�����9�XhcWYQ8L�l ~�K�������$u����6���A�o>�K�� j��7(X�*�7�cUy�pz$ik�~��h�U_��T����~B����{D2 ��+ޛj��= �lNwmv�J���9��Qu�Q��e�	�eDjw����w�-�;6�+�Yk�u�0"<�I�D>`����rF~M���C)u��,���]u���<��[
����R2�L�U_��j�i�~gbp�e|��Y�]�֝`6|K6��/��A�TT��y��,n��
���|� P�.)α����/��Oy��l��`#�`#cP��׏�5t#�`τ^��p�_4m���[^f�Μ�i�i{�wC�>����&&�u�gI��?�J#���nݸmn�%T�@��s������H����Ot{w���<�OO �������&H!�=�˸}e��g.f�æ{4�����>��(�B�D}�����[��9�P7d�X y���/���
+��~냖� ��I����A�e����]̝����0���s�[�3u��У�B_n�]_d����R�l��,D��A�1zQ�9�\\7��cqN�<�O�ap�o�����_�ǻ���g*.�,Ԉ;Ŋ�| �𾈑�^�P��)]��g������Z��6su2.����i���DocK
�(��}��.�� �����@���^+e�o{G^��WaVfC�e^��i
-L!Hhv2lp��r�@>+��(2�I����!����-�!ӡ�I˩��L�Za������h��\�}�sW),֪A��Ș��-<�bR���U�)v�G�hw=s�]��Wt�T������A�~��Tť5���%�Hk��-�<���D��p�
2#�C�l@�5�J}v�z\�@�íY���kP>�����W�����}�v��3z������	0�"�<�"���i&R���ޔ��[&5RAeZ����;�9u	7��9�GF�[�P>+>A�-��sR�5"�_���PuO®Wo[�+]��;e��J�%!ƭ����ҵ�4�����"_���H	�������*�OL����^��&��x�<o�1u�/��}6��9����Ow��52�?���[��jc\<g�c��T )VG�J�B��~i+�ֻ3��{z��3�,��� �(u�Y�-�����F�wN�K�l�Q�m���H��ڂ���
���`���B�+O�Z�y��M��5�(c�D&���5S�t��CX�ӵz�þ�L���\���Y�26�S+M���uܰn�m�'��Xt{�����7��V6���:�Ţ���neo�����,��/j���ک}���>c[�ݴ�}�mE7v��'V��E��߹��*]8s�yI���]8����LsFS`zN� ��mWĐ��4|u�u�J�;�����-r�I�����CF<Y�qqN:���`��Q&~�)��-�k��h؄���I���yv��aL��T#�wh��ja������fY��C�>�)�XL�u���{A���:SA��ݖ��敜�=�;o{¯d�ߒs�]�kF~>������Mm��L'�3����,�:^�ZvU�5���-����PE
F9�-��|H���i�]���.��A�$�*�ete_EEt[<D�Yi
#]��}�	���T��}|LS�V3�ON�O�e9)˂���3��=hv';G�}J�imΝ\�<8J��]�~7��Ott��ʉ`W���I���g��Ԛ3v���ݳ��=F����AyH�ͺJ���_�tPqw���[��x%FȌ��aWG����:��?|{���ǉKrI0�����?��Xfv��
ל�K����v��<&�9�c2�0��M�17��	q�5o��$ i����x(���V�X��TS�1�퀟-��y�鋖��^��PI4C_�]���S�����Y���I�ia�gn�5%R��{�Xf~>�	�g74�~LMy��ven����V��� S%_4���)O�j�r
�Wv3�H��c-�����Z~D�{x������N"�6��OM�`��l��I�e��">���I|�՜�}_�y����s�f�nc-iTQ�w�T��U@�2l7m~��U�SA��5l��=��7x̬���Ύ�	c��G_Alș����A,{������Э:���|�Q�K׹C�]	���X ������ph�J�= ����Y�'�7��`�A���L�>Sģaj�����d*()y��Y�X�ucn��|�־��9���K|���N��.���{��4!lm�')��K�r��4�.�j�oi�!/����}G��Z��IG�q�_�x�M�*�/�#@��R��M��ח8��_(_f鎛���#Տ��4ݰӁ�@�*<-�+9z&�N�D0�0[=���ЁCY��s�oMenb݀䜓.����Ǻ%Q�ĥM��$���H�:J@(a-��D�ʺ�� ����ݢp�z��dVs�bhO�{���x��r;����z��}n��Y��ݕ���霫��b:��k����&���8og�������~���z6d�?,!��t�� 5�*���*��X�=$�a��c��O?����)��W� Nz��|���[*�kf��ao]wAڟ����hW�w��4G��ץ����������Mi��x�4t��Ȫ��a�Ks)�����ebG'�:U�_�ퟗ�*_���n?��u1��Y����[s��=��d��e��GG
�뺃2ޒ>�l�M/WE�����q ��uͷbt�<񝉉2�^w�V٩��I�E����'��S��� �M�x���_v=<�EK�����_�O��P���_#�|�=}k���]C�7���ux�S��g����S�M�x8x>ms�%4��F���k*��Y4�}��H�AP�v��O��v��~F0�(��3�{e��7��m��f��wW��'ؑ�`�!Jn�gzI���2� �Ybcz��W�|A�х�4��=�����
cH�.�?X�n���!��ۻ���Y�tٺxж38W�C�R�uKhI����x��uKe����o+�z&�3��� �+HďI]��D^�PR��[�� oP���٦^�0I���<-�]��������-8�3�`��� g2��Ot���/�#�(����x�Ľ_F\�wFʳ\����Nl�1N�s%������V�"�r�n=V�{���{�Xw0��X��T�b*������|��EN�_�A�D�?녰|]Qz*>����'?���]�:G@����7y��6C�����a=4Cv��Tj�?k��y41�?;܋���m��<�ޱ��}zc�Q+g���{�Y������|�����B����W���a��@�Y#�_¢����0�r�dAh��i�����C��Hr$�~��DHJ��S����	qA�	�Y�8Wc��Q�,|��y٠Ox�7	�����:vnB��s73J��7��pZ2JM
ċ����3��*��NH�2?ϵwZ�³묓��!XE�7c��1���\{X��,�'QC���8&ޮk�;�z4 x.3fw�&vK��4����86�0�Yҥ�)�0�	������_��ڋa��ǟx�1&��G��	�\��0k���#nq������׵�ʵ�գS4��˗���g�'[7k��8�XF�B�7��G������i/�P�ƪ7zE�j�X�7�_ �d�[=�����&��J�^P�(k6'������ņv+A�OH�Z��C����i��<"g��R��v�SO�WRQ���&6�.t֞��I<5�O�X3<��h�-���Pǉ��4���;K�Ӻ��U�����cSk~e9�����H���AI�B�E��]$�VU��[���������Uż����y1�)=�m�����ݳm�j<��<5�2M�?<�� ���7�ߢFrϓ[����(�'�җ�q�ߦ �A�뺆jQ(pΈު*{8q;��H�^��$�:�q>���8v�sJL���
ZxW��?�[��H��@��f?���NB�T��+ƛdP�
 �d@�����{G��P�)؞�f�z�u��?_k��t��o��6x��P �v��,��ފԇC=�����)��RB�r��P��G�.��Kś吞��{è
��ph�v�f�O�\����@�*�g��c���`�4 ���]+�3pi\�#TW�[�w&_�� �5��H��؇x�=�H��;DiM%Ep��l�b��4�3u���w؍�j�سН~�]/:��:�t�ǒ&u�>Φ�NR��T���c{�\�?��	f>�D������jΚ����CB*��D��M����|Q|���.�'��'��ӤQ�m�)q�����G��l��'�UJΗ՜4�tu�h(^b{�����|�J�@��B�j����ZW�oZ �<J��O�z�<#����;����;
b�CI4�F@��t/O`��ˣ<]�Pah��r%�t�qA��Drz_0LP7.����u�ۺ����ӣl�@{ʚHmw�6m�����yS\��:��:3��v��b���}i�dѯ8��)7T�3�v�!y:j��"voZ�l>��^3�?�W��c�J�^$�D\[�{�ך��t���Ї��d��8m�ݳ�J�mn��1���%�����w|]y:EN��Hn�p�W�������4'��?rO��vCW��ݕ��E�8T���g����T�3����y5�?7�94��iݘ���L��*׮��x9x�ux��S�9��R��F��(����CD}
��2J(��*��,��Qq9�,���&�a��G�|*%N�+�P��s��;��EŗD��L�IW������"��o`�u��U��!p<�zn[
 ��
�~�I1�\*�?�f	��H�f-�`��ܞ\��i��T<>w����c~��hK�q(�Q�BS��_���5`��z�,��~�]`��%c�,M>��:lb�y�X!����V��@��r;�V3)� ��&����?�����ުM��� �5pRԡ �X|��B%�e6�]�d^�'9=�R7_ޜ��ѫ��y,�OY�\4]s*���] ���ksR:�k��e�b[v=7��)K�$)(؎,�;ׂ��+JA�P|wZcg/4b����T:?z��O;ֳ#̊N��S7{t�zrm��Ә1q��tu,a#��VPܑz���C>�zn��@���} Y��˛��f��R�J2�yֵzXc���7�
�c("�A��p������ƽ��<<4�LXq~5��j-� �g�)5�m��8���L��k�C��x5�K
�'�C� T�v�=c�^>�����=��`}=7�%�a-�#,��bR�epJ�%�^�-_K�����
'#�v�������_�Òk4Yб�t�ܒSCJ$!��u�mAA�������(��r/��k=EA,dWg+��Ȱ��8�wv��s��-�#�a��ypw��O�>}�74��$���5���j�!�Ҕ 7�'�����Z���w���l��t���������U�qQ97� O���(n���𶒢WP��{��"膔��9���8��5��y}~5�W�ihB%�����G4��@u�j�0���z�r_�lѫ+��ܗ"�����m�8�����<;^���E!~�f/���^�z5�:a�IA�����-\\�IH�X�{h�_���z�h����[a�PU!�|/�3[�̝��oN��27��c��qx}}����2�B�7%�ޞ؀�$�t,C����]��q��n�5Յ6�,��������F�2��ſ�^͢�`%�_�B�����),���L�S�~]N����(p�t�^l ��k�B�R]�9�Q�ڇ�kk�_����q��ރ���駰�D�ŏ�ɜ���C5����o@0�$����z�X�4����cn!��R�lrjj�R��E=�Sq�$g��\��5\�Ƴ���7$�~1I~'\k{#A�kA�?�z�9S���#{{��4��p�vYq�A�w�1dQ��oN~�����a���\�>K���+)�����F;�>ˏ�joX��A�T>F����ܙn����2sTP��)¥�7��x�Gd��'){{�qb5���DD+��s�g3ܩ�\�j4�����~�삷���VZV步����_��]�����Є�C�3�J:�ZXוb/�'�B�i��t�ae�]w��l,�? �԰��J���4�Hl����[?�%.P�uy��G����9�s����y��*�a��:��){{�I��{RF,]ȷ/`�Fս �oC7�B�{�X]�sR���m��nt���Q(.QI�*+��g�]�nW��_�kء����50�����B\����7@�:���U'��1/��Ć4U�p'	`'{��f�,
pw}�p"T��[W�Ռ�_��
e�u��dv��\�.,�q�R\��u�j
'��!�:�R�4Z�ȁd��xp�I���p�s��咏�[���^��C�+����Ce�U��/E5��۟�B%�q���i�_*Ƌ�`�2�������#�T��Ri8"g=�ק{��FjO]k���J�{�-�o
�YY�)Ӻ�M���!���uh	�Yw�w�R�
�%ǋ���z��0���$B�V�{��������P�I��
������3C#��(J4�L �~��E��S\l'��t5E���݃a���p��h.Lu����M����P�7�^uDI��؟�Ǩ�� ]��l�6��.,l*���<�R[��*Q��FC�����=�"��m�;�.�#x ���P� s�۫�~U/��d�sZ�@�9b������Ъ\Be!�/�E�j��@F�Y
bG�G U���6�Oſ�Z�z#�я�La��S���e5���Ԓ��!?x��g���-�1��9�dhC��9�G(˥[6WS�<<�PO�ԲC�P�_�Ws<�G���/������D$B	Ov
YK�Ȟ��eߗ�����IO��I�o)����!4c�:�|�{���������>���y�׹���w��[����������;A��$h�B4����tsB�߲�̧�gZ]�h��������<��d)���Mh����;� ��k�>�����L����oϛ�m@�Ʈ��À5 F ���Է���S�4oR��D�����s�����&3?_�~�<i�Zd�d����&�%�E�b�n���2iD޷x��. ���k��q���۷N��%��ѭ��ss̓�z��Ɓ��<��,�v����o�k��5�ZPj+�IZ�r%�����ٿ���n(<r���G0���B$����x�ld���4�r��%�����������Y-����m��M@#�m}}�g��G��bmu���Z(({������k0_�HCn���C�g�5�&�>qk�S�����vv�2��\wr����ٜ�2��uX^��]����U�����x�����j���	h	��__��?;�I2ˈ�ό虔h���A/�n�ĭ�'�mssA��,B��G����x�m��E� 3x'w��D�5��וLb���`��c�D��� �;
��p�ϟĽ�k�]s͗#@����{�qS�G>�~f�σ�"�3a��io؁R4n�3q�x��N ���O�{������iw��s���t�͟S�t������rD��ȱ錄�����Ԍ,�W?��Z2� 朏8>1��۬���r�_��>V�k�3d*�k�'��߶m�)7�e���%���#�Ǻ>Ǟ�y����I���'��tR���	ٔ��R3����B3v�Ԝ $Q�	NNW�У���[�-/-5S��U�6��)s������תƺ6h�Q"hɺ	�6����Fo�\����	�5�:Oh�04R��8⬉3)߷>�D��\��c��)0���W�-�>8�zY{���Ұ|=ߺ�����_��V�=�����Z��UHA2�q̀���(��3�v�'o���6�=�R�V�d����Fp�eGh�F0b����%j~ V�B9��{^�@�*��"�vj��K�G}V��Au�(m��G5.��}���/��!#��.Tj�P�EeJ
�KG�<ƯDd�G�]Cb\7 ֕�,JHX�K`����9ڈ|C{����ÐO�;Mc�'Ҷ����\��i+ȣ���q�Abx>-b�Ǘ�d�70#C�`��	Bs[�O�yxd$0�41����F�/�4���n-��]A�	��X�WD�,�� {<�9�FH��.��-d�<��H�i| �s܁&tS^�&���H��cQ�	�?(�	��RoT�</W�XJc�"���M�H��&��Pu�;����WA5��	��oej3P�E&�^��0{�[�U�N�K�'a��nGD� �% <I���?��_b��p2jl��^/��K����sZڑ;��I@_o����x1�h�ޞ��FO0Ϫ��--�o'�
�����'�+D�pqb�Т�..
4�
��MH�T0�V�^�K��?KK��*���lM��,�%�`b%�=���ڍZ5(7���m�О9��P�ƍv�#f!������g���N���%���l���p���FM��0��>� ����o�t`�y�߫{�>��*{��m��@��� `�U"�{D����-<��n���3�Zg�h��8��f��J7p���<�n��Jɛ7���-�@����_�M��-P���px�����#	�@�d��11-��G@��|��Ex5���@+Aˡ{i�0����(�8F̗����˜kk����2ww�\��	5Dہ���������%�f�`�� �jڠ��ۢ��F_tzz�2�a�:�C-Ƌ��O�>]�f7��?Uu�_.4��d��E�Z�SPY`�N�^��I��Y��
�����Wϭ�[]�Ե��!�D�S~��e��֕��&/��T�P7�U���t7�+�ra���P��4�5�8O�u��hnֽ&��\p��>��76���y3[��||����n9SN�����✮� �������s"���X
PZ�e�0�o >�3�^UWU���%ޑ��\V�)�6�t�UNx��QPd)=c����~��k#���}��p���o��_��<x7$+�$�m߇��x��Xҡ��ru�f���H�oB����˪�+A�=�ba������P��	�$���9W-> ?��2=�`4���>5�HEZ�������W�LY�+��j~�RX}z�b�X�F	��0-��L�d�HIPQ	:/�&w39�\���q��wL�@�hyʌ@Ӭ�V�I)u�ַ��(� �����U2��fܖ.yg[�7�8�̸Z�r`I��xUU^To�铓z6	��##��3wuL���a7���Р(4�G��Z3�J���b>����c�nqC�P/�Ƅ"3��*�b(��6X���D��ꅃ��JΊ��d^�e�U[�6�L�l$c�L�w��b���i�T���������xU����C�UU��Y8�%�[�x9+骫�+g������H
����x��*e2�`c] 7a��gh�n?'��]�>��ы �A]1r��s�#������ã�%c�e���L�]�\�k��	�A\_W�-� 9��`e�{6�,���ήO-;5$Ԝ�b��j���:}��3�?�6pE*��c�%hȤq��t@d�"}[��8���=�6�w���a%�s�������{^y�ME��G$IV�63���X�����]�Lrs��IB�≸���g�4�]�W9969`0/Y};؋���\i�%�QA
�����p�dL�ߧܼ�,���Y�Ò~��x^E}����������DW
#EO'�����<-���>1����w�I�j36X3Q)C�rӁ<]����1�}�v.U�L���J���DO��oo���
��(�W��"$f�	Wu�z�uH�1 /3�r��� �@[Q�l?�����I/�[ f�c�>�d�Z�����mb h-}�g�P��`�&�H��EZil�\�A$�hvY�3�<�t�b�}����A;�Ryv���ev�ç�����C���.�F�T�)�9%�=���N\��8��W��:C��Dw��tv����_��(�]v�V�
5.�p�+���r9V;�����:�} �OI���W!ݝ{o��f�����5���B�8��@�ي���遣|Y���J���qA,6�6j��틛��OA�$��j_p|$Ş�,���F����r����j�X�|��K|�S�,�6����w�M�����R��>�� ��w5��*!�!N���M=���l��|p����+���􆧾�E��,Y�@�����YBi]�3QI����~9�G2g�`�4ꕠt�@�KDu��\��������h��$2U\@��c���CH0��E��3�#"r�@j<�!3_Y��q{&��]��"�g���"�б�a�\���$)�	��e'����I��J��~{==ZU`N5+4t�K���_�� 9�Ԟd�~����	��"u]Z��& ���ڔ�j���I�$�1����EP�m��c�Յ�:��-; R�V��K^��t*gln��}��>�Xv�x�����_�b�AV���������N������u��fK��>��ur�EA���&葠(�q���ҋqzVm'��!i�i5A+��;8�N�W�g��ۯA!7���sx�O�>Z�:��Hۡy���q�_���u��{Ig ןIT�}H��qA�?b<E��P����U�~&������gh��9����2O�xA`t�i��=�t.�An2Uu�5�t���:�R==��} r���P��"�b����H'N��Z��4BF��̋]��K��C�f"(B(���%5�ײ����2l~�~�u�L����ϻ����-��B5�m@����������J��ttQ�8v�!aq��
��Р����s�)���t�v|�/�Iz�%�!��.a�W�gJ��:�t ����N�T�J�(XY�83��I�wM�[3���9<�xI��\�)�x@jv$�����=C�k!-ш]�6;�?�(�oh���\O��Q�ǎ��lsS��?��A%�Y�z�
 hј�Ls�)$!� ��M����mon��1^6��,�Bv�|����/���q�(������ɿ��+�I}Bx��۬uH .�D?,��#4Ck 6Ed��x�G�:/��$=&���cQ���jS�R��j��]�b� �.]���(@�뢥.]�[{�6S8&��˽n�p�#�h���R2org'�����G}�m��6Ӗ���*\����?3S�<�� �91����܅��j	��E"	���ym�����=bm��+����V�L�}�*����R

rmU<��\|p�Z����"ĺ��'�1�`�*Xҡ4��i���VQ,}-���fހE�c�c����iy@�L�oԈ���̂�D	�d�Ds����P�}!x#�+�?pn���~�\��ut/�h�ǾM��/"�� ���5�e�v��t!G�@���^B�+����.�@\a�����>�MԐ�qCC���OU&�3Yh1Ȍ�?1�sمf�p<�_�x���D��!Ŭ+q i��]�m�'W�鍘!�?�Ek6�MAT���~�8���~��A��ö��np(Aզ�?778VE��7����f�DCf�ۘ�i�2_�%c0q�R�Ǳ-�lN�<A�8A�0󢢢��� u�'���u�s�<Y��B⨈ӄ)�I[ZM�����>�숑K�d�=�,�;4_��F ?���L�9����[���=TG�6e+�@����WS�It6�����Az�\:�^��Q��Y�ʀ��>i;:Un���:r�у*+!�S����(�|HE����
�+�������������H/��pq���ez����(� fm.�������~U�̌��e��A�6c����$�}�{����r5��}���ˊ���t�>%W�����@p+7��Ƭp�밑Y�^��$�=Ӂ�)��� �3��{����v�b��FD�SdD���;/
y���<
7�����~H��T�B������T����{kOD t�~p�A����Ac;t�쟓{�뚗��I�Vk��E�*�"+�g{y��1uS%��Ǆ� �@�= ��Vh�>�����!��|�q�f�1i7,�t�.gi1�����3j�x����;�O�;=�{kޞe	���*y��M_}��(^���.�*7*�F���a�3H��q�(7P�5rD�/�n뾊Q�����ҭ���,]e��#8�ə����R�{F���V̯��׍@�!Z�_v�2p�=��0�+bϵ���P�V�P���S$���'а�Z�pe�g|�Mm>_�Y�!jHN��`2Y�/E��~�SRO^���>��
לMm�Z�I|a�-j������n�2��݃�Au/�؇	��j� v�Ji����QM�G���q�����F�T'TF�����w����}��xDO~ϫ?Ad|���jD]@�l���ܯ��,i�F�`�a(�-�F����G�gi�uKs�� g<s:�χz���M�T ʆBc����ڙV������2+��X�:������2�`���4���B̤�5������}[�=��M��$���4�(�(��Ie�D�HȆ`�nƹ��[6��b���Y�t䚂O}�?AAr�C9}���<r�N{�^�KT��4�d��u�&�Q+�'�n�+mq���TF>��N2l׬b$9��E�1�~W�l�ڭ%���^M~�:��	U�P�������@|�^�z�*��&���tv83M�+u֯�~F8��k
j�g��RV/���xس����ՖP���)M�g����_&u��u6}֢�@c��0P�c��d!1��>7K�<cJ�*��?=6�Ԃ�M��w�D1t~����".+{;1�@G"> Vn��&4���%�(�!�!�i��=�	{�a�6�y���p�J�肐��>��q���f�����X�+z�Lm�+��(�,���v��5��x('!���quT�8����r���?-�&�����#��&�GԞ\�-qJ�<h�9E}� |T�S��è3|����]¸�t	����h�~�j"�-v^I��F�¬CX=z,��^a��-ѣ��eNG�&��p�n�()�iԈ��#�Ñ>Y����3	��ۛ���IK�嗇2�!����'nfiΩ셌T�%�'�P��.>mo^c��ߎ,�����o����Ȭ������ ��};�[莪*ī]{�rI�u� �����}i��XH^$�*y���g����G��7ծ��j"ʞ�s;��zy��s�Trl�7MF��2�>*
�m�b%�u�T"���U�U��G�����3�� ��?f�]��*g��X+�,�*%���}^)���j�H�鞮�,�|6A��:fF�������|�KR߈cY�xDV\�?�P�A%�k�t$3c��2�އ:{�g;^�����⵷;-K9EC"�P��Q��-%��m
'<d�|G3'� -S�U���ڝ��Po�C���04f�'4�\��s���h�Q����Pm�a��`9�?.*���XW�N/�|(I�hKϵ()�B��Ó$�nT_��S^������Ae�����f���d^t�[��옝��ᜡA� v̬��������j�CL|'>%�ToiBz3U䏴����~�B�9'��ʝXy�p�B͎�O���}jQ��[�vLIQ�T�<�qz`��bZe1�h##�ݾT�L;��p5wrr�M�Ǜ��������$+'%ER_Ŧ>�՝-*������Jݵ+M�"dz!/�52��vWf���C{�C
�n��=�G~]�~��>�`W�T)HkU���o�5�wX�7��;�o!�#������u2����P����k��bRH'��f ��q�x��.���/�B�ն��WK�AnAi��/]�2�w��|�77G��
��'(�|�z�G��ج�k��76�s�{���l)��ɬ���hA�J��Nn#H�\�k����F�O\7��8d�L0s��$�*��� ��\f��^��?v¦2[-��(~�Og�)�tO������X�\�~�"�dD��&8����
P? ���b|�� ��=I֝V��y�l�v�3�鶷ہxq�BII_hp��JM�n��b%A����� ��I�x�	���2�K0�\�	�QTW�H�����\KUU�"V7n'mϭ�=7M���J�κ��e�QudTF��-�	%W��9�*(��֧�O���&1��f_	d��/���d��"��W���,;8��Û	�C�a	M�b3b�+8�$2�9��0�^��-W�
�	�s��t�́�\��#�^��Z
.�.Nc�An�A�L�g���,�n?�!�3�4��H���������Q�ǝ�D9�uKjk�]�M����+f0R���i�#��
H�SQ�~�uA��ghe�t
�3�j�s��g��Ig�l��S�:/T�tu��^sy#	5
3y�x�
q�ix3�ٌ�\IKgܹ�,��ʀ/(5n*���=����jo+���.
>S)l�`�)�WD��W����͜Ø�:C�W�#�M�W����rF�M�=}�ࡔ���-����[�Rf'�d%�$����M�F~[e
v���,~��#�y@NoU&7�J
�?Օ�>�9��䝮p;�y�k�I" R�ab��:E#C��}���q��
���!����ʻ�;��V��<h?ݍL���t8��:Dam jO�?��eekv�Q��å��yͲQ�}'�pJ�p����lX}������j쾿ˈ>:�h���"P�?t=Aj��p�[�]+3�k'�iWa��3<'��^̓?w�	����2 z4�K� 	#��sm��s�s�Z���nV=:�?L6�ܹK�3�l��'(����m�G^�$����C9NLЂ�]�yx����|��+�Ꙥ����{�٤O�:ҧ����U˻0�qf@n�$��OC���)�8(�O\`	��݂oF�V FI����P�㱁I����cGlA튔 (�b�E�p�8���Lyc��P�i[
yk_��$�@�ޤX�:����� �`�Z���J���.���:f&��?_��8�����W��g��b<=���Y�a_�djR�{㷪I4��abYC^�����;9�$£\�q*yok�6�r����_���ҷg]��5.���C���߃U�-�>�-m@��8�$:%��ep�!�*>3<�k_5�VB���C�J��|f��{⹫7$�v.�ٙ ���>��_~��#q���=H������,R����Y+��0�:c%%�kR���"��q&����R��V�ww]�5�K��,KD�LH�[切�e�{��&��`�ݣ5�G��|X
'P����Ư�{���@��Hd���C�R��l�HE��(�F����^��cs3��]�������E�]
Ww*�eS��r^�T������X��~��F(����>7�!���w�����Ak��O{���	����:jc9ˌ2��o��ǡU��O�9�c󺐡�k�	]���'�^^�3c��L}sL?����}v����ڙ�w��ׁ����B��<�����Vh�(�t#�	h�9�.���i���,mjT����������������e�0�����s�`^�6�u��k��.P&Z挄o(]��Xբ��h�:A��v#��v��k�h8�h��7a\y�g$!��Z~��6,R��3_N��;f;�XyGH%�
<����/��ݴ�)C�v��J3aJ�Lh�&�2�k}1SpvD�|>DJ߉X��P|���R��D��V�F���%��	ʨ�A�Y��{H::Yr��L�=��[/9�iv�ۛ0������yr���ӏd� ���K�
8: �(�.�D���z�#�J��@膦�v��}v�=9�����9�"-P�E%������<��V�$�;��ߍ -y@�.�d���XHXH������ѥ/cv����_�h_F,�B(I���Î�Z�I��,~�u�#'p�kХ�����$&�,G���cT��GB�3Kmnp�z:���<7���_]��&��'T(^M�/��k����#����u*�9�PE�����GI�F��`gCCA�ngZ� ���S?j�|��Q�K�.�Qv���g���[�g��Fu5_c걫�t""b�\Ei�:�t�킵�g9����ܐ�[t�8��}��U�>���RR�w�JO��9�x��.�EV��l�xR��m0�a��9ӵ��.z�N)@�w�cJ3���eR��<+l�:�Y�z�2�]�l)Л?�u8>��.#��g���zU3��>�MQ3r�nRi� I��W&�RgHڴf�J�� Z�������OW��Y�H
�����^���?U�	rz�U�Mq4�^M ���l>A����֛ޙv�����O��X-*���kY���Ŗ&uz��6�yA{�)wj�O3�k�!�ÍTң�>��� ����X��םi˰њ��K��Y'zJ��%� ~����o�ƛs�������r�~��t������ � �Ł���/(T\TB ��iuY�۳�����$1΁�_�F���B���L���JU�����	pHx�ZM�޽Xn�<���^��m��4�7i�/k°�� IR�1f�Y��0�?AE���������~���7fU��ɳ�-W9��7=�Q6���8	F�;��xڤ_L���&��`J��������ԓ�F_��Mv���F�S[�U��bi�T�E��0��h�A�aYQOd���@(���H+���Gg��2��5��uYY��,��˃ڒ�dj戴���b��\^�ܽN�����+?��Qk��F&ޓ�\�ذ}��"��an����(�:�O���������/xZC@"�t'V7�NqEE<-�E��O�hu^���ִ��%�z����:�]���󾑹ц�s�r�d��q7�w�DYAO��Y*~��͑l����D6D��5�՟q��M��y�p'�?�2$g�-.贅�(��=��Ͼ�z�	ݹn% 
D�g��]�����T��`�yR��R:��n�m}�_��@��!�B��Y�d��O�����L }�U%��i�)<�a�e��P��l�IՆ~��ڪH�cý�ӳ��js���H���uW���J�s�fSih�����d�'�'V�6�O:=�sѴ��Vn�gOH���S.]Q���ŵc"��\E2�!���P�D
1>T��J�	�7\QQ�tGyz�h�ط�x���IHx����D��<�8�Y;.���m��jY���o�[���Th�NF"��cSg��5� usS�ڛ:&th�cLG����$�-$ޅ��n)fҾ�1�}W�nx���u��oa3�����&Jؼ����qz���q���q��3kNNN�T���pu�ίB�>�'�$��t�zh�G���R�:�X� ����Zm�ԝI�ߢ��t�9�87����m-��CC�=Q��' �W�<c�8v�wC�-����C��]i=�!+{�E���G��PgC"���Y9k����ኃ����[1��Wĺw�����5`���Au+�����@o��UU�ɛ�roS]gZ3��(�p%:'^(yCG2;A�kT�W]���1���v��g"�ZZ��M��4G���u���O����gĭ��Bѥ�{�p����|T닢�4�'����i6�a:El�N6Vإ�~4�/b�\��}*(��朚��r�'���^�}T:;m���u�Y'�dF���Շ�A�K�k�%1zz���:����B�H�6	j�.u�8�g�/B6���<�_�	Ci�]�	yVp5y	1��$_V6Ԫ����.#-�{�r����p����b��*�7޳�)f��[������.Ǫ�t ����vA�Y=0y/OZ��YR�/q�M�u��;�ݧ�ٴ�#=c� �
(�Z�d*w���"�6}��Ɔ8���y�V���B�f]��S�jlj7J��!�c��kލ�b-B1=��(��@�t��p���n�R�´�9)Պ�����K�V������!���̀5ǰ�m�i�g7D\"���L���{��B�-����[^�����ٕ%B.�xS	�fݚg�;/K��K��6��&ZZ��A�2����&I��c�6ixkP��z��MW��2<D�E����r?���e2gj���� sQ��`J?��	�������==��G�a�'�d�1
����g�	���XHz���,�6��!LK��{��=&��3�{g~]��n���ր��޹��_��"w���hWE\��V����o�:�Zh������l8|��@
�J��P�	$�S����p�TTe.�.s�34;�Q}����-%"�����K���XB���fF���V�a5���r�lN}]4�R��5��gE�!�'�%C/͌:&g��_��x�{B�DE��5<eWh�$�-�6%��u'��V�E˝�i�ˎ_���W�j�3]K0s����D-o{��'�bz�>�N�@j\��ZB&J'��D���g�G�~���FY8j�<�)ФT�`+j�R��"ٝ9�����Ǧ=��[I6{3��;������I�l���Xj9ȝ s���ތf4�T>���?���c��I��^x�|��q:�
���� (	�W&l@3������h�,���mE��Le��K<�!?wN JL�@����t�Zg+���'p �*4c�<��-c>��O��"�[<�9��%`��h��Vn4�0Q=A�Y2����$�-_W:X���յ�{\4K���/֨.�M9$�g�G�gK�a��I���<4j{�m���a&�l�����C���p���~]q����|;i��ى&ݹ�\�i��M#�x�����~t*~<aI�B�s��5K��A���o<�%LL��%�����W�4�wD����E5��)Y�i�j��������vHl�>f��=��b\G�<�Q�e`�Emy�r{{��@妫W��G�G���"�@G�:��h�Y�"�&F�Cw�fI˥�վ��c�؃�
�;���Ƥ��M�����u�%�nyU�YA'X¦_R=�Q�E˩[5��g�b��5[�[�F?�h���=�X6�y7SR�;���I"�M����7�Ӎ����M'�xjgO,r.��s_�[cS�z݊�c�������E>V_��X����`Ե"w��c@=�loV���Pxv�خ�Ţ��-�n���	���^V���/�䓿ہ}�󳵍XD��T��ms��2�n���
���✖�If��uta��^f����`��?�^xTq����y2ZT�ΰ@��qѕ^����/�E��]�g�,�3�Y�vCٮ�Y���t�=�y�Y�qt�Iٯ�g'��&��9o����l��_T��)V�RhJ��4���n���H�L-�G)27s�ǳ:I��Y��I5?�YR�X�F��\v���;�S�m���k˽�����;9�C���7i�]���8歕)�w
	����]u�V5z��`���	BB��}j��Rô��+f�~@j���a�0�!�N�g�4Zv̤
�B1]���$,���f�����e����ە��XD@��]?�e����綪H���3x���q�/�.��)_m����͎-��yx���,�(��1s�Ǎ:+�C���K�O�Z�W$�F�*/�y�.�b�)Ø�2��f����Sa:����F?���q�G~��D��9>�t�M4�v���{���#r�	�U똩�c�ʫht�g�u1�x/����es�h4��L�?T�{tnt���v��W�%Q,��vo�N/Ifv���{f��;L��fVE���G�/��#�.����"�[b��'Zj��?R�\��_�c���U�* yKmj�|^h���L���U��I�&P��̊�}�7z!)i����Ì(���s�Z�z���7��uUڽ�o�3+ҿ�&�o��j�|×��b����V�u��#�������&D��nX���(����_�����v��jm/����LN�n�m[p�bnqzǏca�! ޅ鑹��%���������h�5��E�������$�Zw�Cَ�/�uh�qU����w�2�p�Xտ�����k�Ӳ>���3ή�t��IО����W�wwcS�,ރa`��dㅫ�j8������[˅�鞆0�R2r���Jע�x� ���x���s�+|�����a
�M��/�.z�ݢr�G�
:ť_Z��jǡ�eǼD���%k�WR�XL��f���)��e?��v�aXN�mM����-4'gM�L.���f���m�4"x�z������
�g<���vy.��E&v���{�X�o�"�
���0�SJ�]f�:3�8�[��%�6k&�9�Qa�|��kc�VK%�� M�_�0�y-7��CW�Y��)�M��w�����#*X)1���x(t�dЈlʉ�~��]���)y���Һ�3���wʷA���v��=g��[A���abڌL�F-k:��-~�Vqyy�9V05�Z>�:l�oG��Ȯ�f��h�O��=�n��S��R\���?e�;n�&>K���v��(�`IE���_���i�=��'*j��9��d�p�
��Y��.�ԯ��+�Soe�)�S����.A�>�:�p�Z�����5웳�ޡ"���έ�'-��蕷�rI U�O�{�*�������e�������+����\�v5Z[Ӟ=�My+�E�se����4ߵ$�?eEభ�1��
KI6��;C�睎��YF�=ȜBjZ�� ���~��
 �Ȫ��#̱�/�E��r8k��`G$Ѵ^(���:���TI0���F$�pa��b��]&GDd�$�x�����<�OMnw���{�^���z�sjΟ58y39�>�!22s����W`�+��b)��v?����X�a������e�������|�zVs��A���!�s�o��v\L�g�	������2 �,ƃ�l���š�����;��	����t���۞c��7Y� 'v��ΕK�R�7Qҷ�w��Z�I�<O�mɰT�M={WW��Ee��a�[�K_��b�>��y��DAH�<e��y�:�&=#��K�2��OJ��s>M�ϙ�.�x���9��P���s�#�; q�1,����KP���㷦إ�,�Ym� ��+ ����M`*6}N����԰{N�[2��;¹jtQ�f�-����}�B�[2F��V�h���2At���gl��;׍~m�Yu�+�2�	���K!W`H�[_6��EVk�Yb!���D������g��;�[��.����q9�n���(�H����B��A^�����I��=l/�D��^��h�cQM(�_ZcbQ�;���CٌOm׻�5N�'J�lm#��]�B��f	������4�`"@�#��o��8j����}�x������Y�W����,y���|�66��J{h��Y$���$�����5�� i���G�e�J�}�l�uk�4W̻�~����O�.�	�n��Aײ���F5[�z~�wo���+"8,t��e�7�_��)������}4�1�ކ�F�A<pP�,.?G�ï��?�8$z0��,u|{�|¾m�OR�^�pFb��(�G���<LM�.������L@� ��?^|d]����n�Կ�����J��1�(��B�o���QN��f����e��T���h�ҳ��E�]�0FP��Da��i	V-J��u�»�k��P�ɛcyN�Yx<Sb2�K@Y�M:�w�n�"!sse?z���l��L�0#�'��n`�� ��G�&����<�������߶&���4�h�<�̊�m��20T95��i��?OH�	�'������}C� ��h�'�s-(��p9(��gM�_@��30N2��͗F?�65GȮ�,��r��3Nb�(�V��7Zs���*�Q�U�F���ICޛs�����c*E�d�$iD�f�A��߭k��N`Ys�X��
�r(`�H)�F��Z�Z������X^^ŝ�&W�sa]Ե�p��T`�I��f�+��v6/��aR���O;bG�%�h�����`K��X��d���h?u�|���4�"�u��+yC�س,��Mx��o̝�}�Ǖ����&�0�)�$���^�ɳv�u�K���.M�D���5}�������gM���[+$��v[/���"�I��h��w]�}g���N]�w2$��@�Zu��P.:�wf3��b}@������D1	���k(QS��s{uOx���p��Դ>{�ë�n\.�����#�"3�#,Z|�i@���x`m�LJ�M�B����kتӳs���m��0X�A��l@0�aD�Į�0�~��0�[��7����Á�2S�i�&:�vmo�i�?3��(��ϹAf]��B�|��-=�dc,�� G��+�*���TJ�53M��Z�9�&B�V'�r$<��ڐo��JRe���M�F���E?O��/fћ!5��fW�������9nP*e�U��"����6;��Ђ�2U`V�Z{�i ��4��g��У�/^� �� �{J��M�y8���^��͗;�B�L��}P�5ڊ�� Ņ.�e�T�2�5ຜ��YJ� 9l��L�de=h�]�����rt��g(4�@���.���4|��ϻb
�ax !�Y]����T؞)K������K_�g6�^�G����4W�6����wA�(��#�)[���g������z�a�M���U�*ӵ�?���Q�AP��|��|�P,�m�s�Ű���'�Vj�l4� �x懟T,#��+F��L��O����^�!1,������ɲ9"Iw�O�����9����Ui��t��@���m���S��k:sOTc7*8��}��v���u�����zi����Q"o9�=4>T蕬b{V���?�ԠP�����q�O��\n2��?w��f���+�-�=����p׭ �~���
/�k��A��ݱ���2�r�ǟp^ԨK{�Sô��8�
D��fX>x�>;{��0b�r2ܡ��`\���5I+莾��������֟4=���L�E[�E'w?�V/�"}�$H�V�؊�O���l~.�a��2VӍ�s����ኗ
E KG�v݆Fge!�n̿,d�,�y��o���ꑋY��k�]S��8����&�xg�W��WCG�v�42�Z��SC�����	
ڱ�d��u�uiN^�]��L�)������ኙ1̠��u�- ��9����,̸M��bb���ݭ��[�ڹ�p�^���������rٿ"JO?�^u�!����|��G�;���.~.7�r��OR�X.*���c[��*�	���?�,�M���wB�g5���Tf���z���sv�����Vπ���H����_����.�gF\f2�.�0pz˨.�|� �z�^:f��Z (��i�E�j����!G-3x��c��9Q[���kz�<�9�Ӿ�З����,'�Gtq=J�S��c|]�����Y ���;��?|�����$��p�cL�ԅ}8Y����I�B�^@S�:(ߥ��E �k��$�۽�{�E>����B��\P��ڑ�D���g�	踄X��%�!�h�2+� ��%��s�� �X�4��ZaUl {ST�,��C����br%[��z�nG�O �[Ԧj�.<B%:�����%�t�ѭ�5K��Ǘ<3�К���,����fE�ui�����"..<9e��[c�4��u^;�ȅ�+{�[7�KH>�QLt�l��lV�+�@/@����+�F�JA����9P��Ũ�֢9�k��d�(����)��i�G�� ��G�9`�Wt~�͓Z�E���H�\��!����~�Y��*�`$���ʡLY��2��[3�u�X�,П+B&<�VG�����O�s�?�����z��1��۳g�f����wb}G�eM���kқy^X�>��Ӣf��(�\{�sy,��6vT+���v?��*)�,?W�h�^�8ُ���$ ��o��-6�2�g��%*�jo��63;Vcv�����w#h),���ؗN��Ɖ���������`�{�9��2�
������OW6H�;N�\ u�tZ�Y������)��j�%��D��u��7,�_S[@ݪ9�`�.g=��=�H��U��k��B�/̊�K���"!���@�M�� �ޛE��-�ܭvl��Z_\HcP Q��R���~�S�-�r�_��Ujm=�.n�/��'����#т��/���������nra�=��z����b�h�@7��ܕG�.Ztb.lV�\��J����܎��~$�l�b�yV�ʎ�Zb:<��~��z!���K���B��y��	��7m:Xس>Oڒw+�ж��J��w��C��E	[SS:�<T-�U�����a��>�X�G�v
�h1�����쇊�"�!k�N�g��N�>RYX�'�W���|;��`>fӯ�p�W!��R��r3���$_��Ix*�X�ey���㉢xV�ݝ��%RO�~��"�&�w��<��gV��=�D��W�/R�:��������vB�|��3���~Pn휋/�a�g�O�a�LN���m�F�)��`Y*�R�ߝ�0�:���{��#��d:*,I���_�uP�n�'�}��f��Cy���+��no+~�'r�z���1ܫ�|$q5�$D}�U���)]��;���:!H��?�^7:e�tV�9�ś&>�$�\��&�2u�4	�R���K����v�7~�ڐ�����6~o�����$�Fp�aU�q���V�i{��;S������*���!u{��[��s;��j�c�d	��f��V�&[5���:� -���ocF��,��
�����}4�K�(X�f���-(�����W��V����57+|��~�U�|3�(��q3F�Ĵ���m[�G�0A�æ�x�����p��rč��;��_:3��t��p_�tj��?�x�+1i�7G��ޔ(��եy՘��?T��#��,i���l�!A#������8��B�o���?Җ_y���X�U�����p}�?��:,��{DAE�E@�AJRQ��.II��4�G�����Jb���$�`�y��<����xyy1g���}��^k�9@�}y7;Q4%��3�\d��{��_N�^���H�B���}YeX���A[�]峐'�|�`�Q�t� ~Om��.wP~���?��אv�T� ��;dږ,rDe���>�CN�A+?�y���si�,��%��n{<�9����%� �z��|�]s4�����ǝE>��a'4�w����@�b����H/�X����w�		��w��G��-�O�CK��9������8�8f��P��G͞���y��8�o����N\���C8!p)�XZ�f�r};��w�$������z�w�R�|�~����)Hv�����"��~[GGg8�pe�G�bz6h��_��q+�mY� �HA���?{�,
nE����;.�U�yrs��9D��U��>���T�Ĥ �,,��֨炵ۺU�}c��	��[<����FW;F��Eo��k�V�����՝��J���B �q��y�|�|S�D$ dθ��^���ɣFw�ݧ#�n�ē`�.����_ 	DO���K`�ɾQ�n�U��.$�|�:>B�d'bE�y��6���� ���m�W��v8���8/��D��]�`�Z�v�ی�:�f�?�6C��Z�YN�����
Џ�s0��s�Ah��}�� ʅ�ȩڋx2�4���홓x���ס"((�����Y����KST���(�� ���)������$��'�}�-�j爇�W�8pؗ�q��FvM�ģ, +�?�"�Lz{����%�漨�]���!Ga���^�D	�WeO��Ou{a��"���*��98t��!HV�exwP�k1�޿�y�~�N��YKE�D�����{b����E0C��r.wb�;�_�z=��o+�����J D�����R��r�
ѯ�Kɔ���,Ѐ�M�,��Fx5d�O��ѯ�zH��������l����R|<�V��+x�����Q�ӧ�������..[K���	��G�Y�@cQ7��2nm�+��ϧ���c��&v�:�����{��9.-�,SM����ҫW��h-�:�N�$;�3(k�������e��*�?�j��WZ7��(uHT�^��P����)�i������э�*=���K��/�rfڢ*���`uwO��)�7q�svW�'w�"'�9�DbwP��5Qk*���%*�$V��l��)f;��9{Jٳb��N�c&���,���I7�+��4s��p�b�cwm��E������)R�YςkJ��w���R�0��Ώֈ�xy]�C�@Z{ըw4n�7�����{����>���xS P8�}/"��wB6=ȇ�2�� )9��e:<����n�?C��\a�)w��� b�x��X���+���C��}��.����h����dw�;̡�F�����v��c��>��Κ�+��T��2�_5Y�:jE������Zj;�Alnr)�^x������[2{}r^e�[���1y��^�%�D#1��p���'�4��o��NI),�I����iHx�̸����6H���2�"���>���c��=S�����j��eW����e��0K.���"�:Wٓ�M���J,���1V�8�l��:�<4�@S`���s7���ZNlPKK��5�3;��!����g��ޗ_l-W�	��e�-�Dॖ�N6,��o|{���d�<�"���k��@r�����ƁCbخ��|�T1&��UN�7T%�Zak��VX�BBO�1��3�x��'����Y b\�@3�()鮑e�����N�Q��Z
��(��jCYWp�R�Oi�����;u�[�	[��$�K����$px:SH^��
U�Jt��{ �@2�Z�Y��3k�~JH��H�_h*#��xm��)���&�7���f����V$�U�
xl��y���WM��+=C��+�����ѸO��cw%��0GNw݀`�w|���|quS��`�'5�E���]vW��ĩ�	�K��̉IT���e��w,O`��,cG�����xKH;�x�W~]����P�}8����p����C�~o^�vnع���5
��2�Z�=ѵ��v����>��}v�1�L����q����sj�!.mΫM���/�S�J�����{U��0Z��g2ҙ�$jf%P/�%VP���O��8+��w��L�MX���8��w�A����aQ������5�C}�wJ����CTbי( �m�����Y�%��e��r���;��F3�$��EA�-�/�E7N@���&�]M(�C�E�"j�X�#��_Q�׆�x�"73Q>�%	���Z9�����sG���Y�1�9�wx�-���w<���-XOXVơa?�w�
1�e��+VA�49O{�#~�J�b�	��>�1��ןg*�������@��g]_�����L`��֔N���(�(�*�'�i<�3?�<�bp�EII��.>I��3���l5S��	œތQ���[fD}U�f��x/|Z�<ۢH�쇈�v�����\WU�2���qy'_Ֆ�Q�O#ݼTf�h;��a&A�x��Z�е�_�W<��h��]�7��&,�o�-�.��g]AA���ݼ��),�m��9c2�9������lP�f�I�y�w+�d�zr����0㗞������=�����Ft$��R�/�DC����Ą���7��jj;�����~g����xcj�7,��r>Np���9ahdc9 k���^xچb{n�c�O䔂N��	�p�ݨ�:bG�MA�bR&�B︗�[�5:�/�)�\�d*Y�'�{`�:F?8��S�P�e��V��V��\/�]#Ǣ�>����/���_��-�bf�����7�"R�I;]����Q
~c2��;���)�t��J�B��]bV��.�(|��<e��2fw�T8b/39� g�Aby��E�a�u\�2v9}8�8�����~��FY5�h�0�w Ȩ��+�A���51���J��ϓt�Z�;p�P_��b"��j���?�1���/��2����:9u����U�?]5��YTFu�mq���x�[��~^Z���X�����J�M�Z��]A��ԲL��5F4���Y��W5�!cq�,rq^�>�������3K�A�χ�jČO�u�\f����t�ݘ�Z�����>���QSY��W���N��գ�Cp!���dC��� *M
�X�P���XeKdP?Z��1P��CQ\�zG�lN���
~�ʯ˧�&�-��=)�m��%� �An=��������˲�w8Me	�����Hs+�o�V��*´�486ۀ70v}��g;fџq�Ӱ����f�)Gwj�`�խz��8R�gh>}S�KC�g�</d�
;S�����䯏��e+��'"��R�����,�e�bK�v�-PU���:�I���V�i���i��n� ���J��K�}�����\O��9�Y�^8l=`|&���_%�]��j��v�\�o�s�F#&�����0�g��@�����}=��w`�R�S�p��� ����?b��Io�])���Z�N�׊���`���sr��}
'yg�;�ٸ�\ʅ�.�
{W�Ϫx�H��07�v��%G�w����]��@"�R���+6�S4���\�<X��<PռB��N�TV�Jp�$�$=�P_?�q�9mɷ�N��}�����q$`.����un�}UG$�sGSՠ7O��A$y+^�K���\�~�|K��_��9��>M�:{���͂Ad��M��2O����Y\�������5�$��АW�/K���w�J��3��{�l��*4A{�|����^fS\��ɳuȬD��&���0��^����Y���M�	�Zf�������,g
Ҹid�;u,��'M~�p\a���D��v�!��k�X�9j'����D||Ӎ��x���Sq\�1G4�尠�Gʘq�mX�q�Cx�+�s֨�^lR�<3��Ь�<Eqݝ���҆�~U
g��]k$+�#p�o��=ӼW�&�R5va�!/򉰌C&�↯������B�~�ă��;�`0����GyEu�
��6�`Wt�2���Ts�6�v'��=����ә@�"c�w��쌺Ys*%�)A�L���!�7�0b�z��-�-2x���W���Xe�0ԉ�Ɉc�}��z?���G}w%%
{��/R�A��9� %:��j�����M��g��Q\)R�Mb�ų�]�aY�qT!��Ƅ�2<"W
q����%�WM����8��j�8��UvÛ�DA���*/���	�XA�홣h�z��Ԟ5n����ƔI��ry��<�i .μ�|���}֫0 ��I(���!b�<s����J��`���(�ӿ>U}a<j+1�s$$��#��Ӻ,4��߅}�[аע}��f�`��s}�6��;��M�3��$<�Б >�OQ_�y�Zԏl{��{�z�����
��9}9v��%+M$���p���E/����N��N��kL�C��H�Гn<cX�\���/�L�����O�Y8�pA�X�wp��~H-���\����pض,q�/'A�:�����V��5��:O�u�vG��8b�綦6{����R���w5I��<����l�j�ɧg�R��P~8����V����/e��t���w3p5u�@�g�ӡ�9�@,{��>.�I�����;{����"�Z�?��/s��@('���K�h �8w�K��)�-�`�uw8���"^	e[%~�W���q�(��\i�	�J�L}O�34�oPk{�;oࢴ��zN���We-����Т��S���%�¡�{)΅�ӧ�45�֩�҇�@��'�����]0�{-f}���>�:��}y��5i3�<O����a���rx:0���w׏��D���I��<�o��-��ځ*�lo��0����� ijz}��(�R�ng��d����$f�(���浑gf���;ļ��	+1�_=X��8Jb~���/Sf+Z��-z%�(�~,��ܓ�n��V��y��N�:�"���K����vW�C86#ޜ�a����`d��f�o̵��X34�g�JM��<�=1:��<��'"��jC��.����6�;[kyu���A5T�&�f��3K�$�:�<���~ؓ�a����F0�v�����)��~K�SV]k��@��s�: �'��qB�L��R�)�eII���נ�vKbȏ3!Rqhqw��sU��^����ZyI�\�k��,w���s}�v��5^ޛ+�Z}��q$
l�FL�U������
�sP�5w� �@ �fd��Uc��0O�/���Yh`�1����b'�n���=Ą�_2ߎ.�ogbFy���k��k����F�p+U��qy��m��m5v�=[S.U�%w���g�4��㋪v�P���}V����A��l��y��q|�}� �~����)fq�&)��?bbV��H�)*�v�	$Qp�yRC�k>,��q�ȴ�CnH�t�D�袡-�ӫ�Wi=�3U��$<}�'�J7dO��s:����T��j��� ����>81+����i��S\O6�;�BBE���3��g�C��ߒ����։<�{M%���*�@���O�6�E��|�Xp�z�i��4��x^��T���43ZZs1�}lD�>�K��~#��)�%v)�W�j�㇘`�
�TX���1�c����G���}wR��wܷ���ǄF�ϷX����r	l�8Ծ���78`�A�柚�i\�,wAW�vKH��M���͐��B}�.v�c�ԙ��7�+_����s��@�=	n=�d ����.y�V$�ׯ:�S�L���=6�N+Z�A�󘔔%���%[ِ��ND�,�(��f^���bgC�}|��W�<<$@>>�sU�Z�A�z���F��c-9�9d��m~g�^������Ξ���e6�s��}��0��EF�Y%�a*�� Y̛�{�rE-sn�{J+EI���k�AH��&�F(8�Dr�I�YX��ry��h_��k|5�ס����ָv�_��9̲̔?ix��]w��Ꮾ��K�^�A�ё�l���b�ui�'}�c�ʲ�������,y��A��������w`\�<`ld�G���NJA���7B�5^����Cc��([�޷�458}����:)-k��`��qGb]8�ɻ�2�6�5��
u��]�|�-T9M�w�m����^mT�ij�L.w��W}=��(3�@�X&k�hZ�Ϳk�og��4))(�(>`�&�z��Vj>C�x��~؛�5�a��\�d=/
2=�ʳ��ۆu9gS��\��R�z<�3ē0:{K����R��X�e�$
��>��Ii��b��X�_�0���Jӛ��{25##ug��4=�?:�XgG|�Av�kp�Khjn)�/�/������D��*Z��F��H3+��6�^��]�ޢ��%{u�%�l�%myM��c��K�h����w�C�����^�m��r�I|q��f�7�
�r�~F���;wB)|6z��-`KfS��õ��ʒy�n+s�����.^QZd��춓E�Y��WT��G�h��r\z��h�_1
@A-��އSW�\/ }������	2_�e�Tfi����n2���v�b)�Îu;u��.����r��v���Aibۻ�=�t�}�P���ۯU�K'�|m�)�:n�q�ʬi��Q�P3��R�I�7o����E��a��-���2VG�������q�)3��$��F�b���J��5̐��UTvTV8�Ȟ�:8���П��7��=�|�C�տK�,���X�k%��5�X\Y�y��;uqN۞��Sx&�+p��o��Lo�0lMLJ�` �ԘvǑ����`H�_�ў�f(ΰ���#��x�ksV>$d�ͽ㞰��JQV��#Z6�C_T_�|�  �T:H'mpl�m�]��u���Qѕ���C=�g�6����}�3i߻Uֽ� ��^�w�d��B����$��x\^���v4��26��_;qfk1��ˇ�7��W��t���,�gZ���ΕTf$�r�V8�ĔHoo@�/�-]�FS$1���#��.�a�/N-t���ר�_gnn����`1�{XB�{�H��cԡɤ6��
z�e`Э�bt���4|�#>��&��M��ZR���#�$5��Z���YB���A���b�7d!��^P����pe�`��m`o���ߊ��;Il��N���Գ�����ڗ���öRQ
�^x*���fb=���Ԝd@JT��	��#A��c�as�X��QzWG��v%���z��d��U�ڟh�H�|��h�M:�L[V������_珗{�o}+���BL�YS�_�̙��.�F�!S����N\���@,FD��K��{e%�&+�be�q�[��2mS��Qx:�)��Y"�@�D��k���-[�|�"�C����4��C�AC�)�[��<Ej���������	�,22[n|�
���)��[*/ {��O��MA�pm�e-��q[b1w�z��P��k����!�y�^[JZ�&e�l84`$�@����|z�~N�IH���.�w:�Ƃ
�;��JA'��ꩃ\���)���"g��<�ge�x�&�ֽ��&�D&�./��o�6��E^������gM�8���hA*��Q���͑r.�G�6b*	�
�X�$b�RC�<��#��B�W�]��N .T����xM��fߦ�c��J�:V���:띞���M��(�$�m�C�^�{Bi�I���>��q���7oj��*�;�vwo��^�h���6���v�Pt:��x��1��W���AQ�b�@�[n�C�^M���Ҿjj�4��d����^u�6:�8�E4+�����N��Ó/G�1�gUC�bbp?�e8��R��~�J����#�T�sv���Af�Hsy�{�>��Z���������}���o�[O�{�Bng�@��ᔡ߅q����?ȉY�+��B{3�����7J2?ɚz�����M�>r���׫̭���U���RD��kl�˭��'�XU�UWΫv+x|~$)�VOl9��R��Sw[��]�S �Z��XϥãI��n���"�;�U�P{�
'' ��M$��7_`�(�Փ��M/�;3%�eq�c����}x��j�A��p��ҏ��X���م�R0����P��.y��w!ZL�\�9IM�#M٫�7y���\�����N��YZpK\�����4%Z��>"�DrI�|yW�� �i�a�ŶNV��;:���է�
�a8Vi'b�QY�^Y���(I���lLW�9z�X�Ծ��r�ۣ��3xѴBP���JK��+f���5]�c�v�ݑ�]���W�F����R�X�%�0"�M:)vv�����#"�6��*vm���N�����ط�x|x�>�W��싦����/���9�+�����g<e�8ȂG��,��	����X!l������� �e�ݜ.a��NQe��s�����6&e�u� ;����A�{>�� H�=�֧������K�A��-#b0\';}��g�8<������p�*�;��O_��kW�K� ���7=r}N�EM��51��L��NYD�<+�|�.� ��V�J���>��0�:���R��1��ۓle��X���hkda�b|T��[�Pw�M�?�������xqj� B�cH�/ՠR��ZsߌYR�g,�斖�������ɑ�#����J.��҅w��
�����֞nJW�u��\׽�(A���½pF=G$#��D�����.Wt)[�aW
w�~��(ߜx����{T_iڮT؎�_�y���J�F�����|C����Q+}��
�ز}v��<��[�KK1�4}rvI���cC{��O�dq�C�>�h������V�xEݘ�|������#���('�P%�`WEUo2�p��Q�䴍U�/N:Npb�@�
sԻʭ���4��	��&/ ������ߋ��������t7��$��(G���W7��yH��x#�q"pKe"�%��'j5_��ks�'���D<6	}L�:.`�GP��5��.JJy@C��ᖤ�O����� �<5#�ظ�k�Z��5��Z���2[���d�DWyW�U���;�;QR���x��^�`�(�l��^��d�ڟ%���Y�@��რ˴��@Ա�Y�ch�tJ�x�R�R7zrjs������u���K��q�N�\i۱nq�S�(a�d�i]���4��Cv�?ޮY��bd8�L
Q����Ȃ�Ȯ������_%�ϝ�/�Q�\f��{�
�U��՞*y��f��a�6�@F%������U�D1os�+���R��E=��{�G9���+�lA5�z�ѱ�D���)Xtl�+xCQ�h|؝̹>f�Ha�O`��(/��Zg�66GZ%�&���~��
M`
Bed�b����MΔ�a����`qA �g+*�-�ndx�_~�����.3e���;o�������k2����p�	��>�2P�9V)�����-	��O,������Sz��i}�P|���ze��[wY4��mg7�C(�J���{�3�- C(a@qʫg�����;���3�V�N�*����Z���_tn�^e��'��~�����@ӥ"����ROv���Mi�g��#�����
jNO�����l�����b���7" AB����m����P0�(1|ېK��Rc{���a?�kܙ��t�_7�_5.�'���"�1!>>Z�N��"����G���+�<�[v���
��.����ևd]����+���	�Y~Xz�F|��S�Y���;�k�]45�qC�O��a3Ϗxy����dd��t��Ź�����L������ԅ|Gu����B'6W��.��j���t��h�i��a�U�����r��McuMs
u- jt����Ԍ�x@�y_'��;��YM0OO.������Q1c���E�V�>�? Қ3{8�"�8����L�ݿ0�J� ����HF�D�}�A�"�L��,������bQx�NO5m��?��q��x��ho]�;������ ���`����i�f�GwK��O�uV����ڲ}^ъZ�>2��W��Hu�`j����?�������uU&u���u�cBB	v�	��s�^ɜ*��!�y��b����#�ü5��ޠ����W}49j�It>��$ޟ�4����	Go�\��t����~���P���0n�|�n�*����Qp�٭�Ƒ˺��=�1�&Y��{�	k-�X�����H�o�-�e���diHAD�9^�8;O��һ�W�3y��*Pc9��iN�&NN^��.�'쾉�Xp�r�yK�'�S�_�n�:L��P!��#�(%w4�)jf����҉����Lz�d%Έ�6KT����y��I��A�௓]��NF��?T�)���o��bwM�	eXc3D�v?kc��������	�xpQ�||�� k�4H��h���{���I��Pcr��C��tֶV��n�=�W.��8,H@O�;�z�#�F��'}��@�dM{֧O 8�ө}��GB��|��*5�iI�u�B+K�ЦW��T�֐��d��)�i@��u����ǽ{�%���XL��;V}���OuI4#|f�b���G�T�7<���`������+��#�N�x)�������1�B����".����Zy�6�/Ga8�؟�f���f
�-�E�0�o�<R�w��ɝ��u����C������S%BUmJ`ؼs�X/Ǹ�<�verw�9��-H�P�|Ҋ��M�/@�S�{|�(@~�I�m�QI�M���Hy2�¨n���ʠ���(����E����'�*$����c�"�G�tw����e6C�%v)�oޔqj=���>p3����hJ�B�T�qH�� �����w2QX0~B�ˋ���j(�LJ�&��xE�i1OE)�;XG�i��C�_�H���5���%7߅�|D&� �jʜ�s�V�s1.2��#�O��l��:Y��#)X�ۏ����^�l�7 ܵ�����	�ZKsL��("��+|�t���e7�=^������L��z>��<���&����+��Nzk.;�e�:�^=�^I�˩5� >��4(O��{5���7��{%r�<EP��U��3o3��~��+��h.+�r
"��e	5�|
��5*҉��O;�Y�,ߓ��z�o���|Vjd�����o_�пc�^��,O��75��"`n��gz[�N��Q.{�@Z�Ίԍ=,b2��2��9CD�m�s���ط�˙���Ͻ��{��뵡���O��"�j�?����|F���Z�]�Vj|G8}�C�?�y�~0�����urpȣ�<��=Gz�Ma�r��ɚ� �4.a��&�C�_e���e/󱐌�_��,*�ɷ��Fx�F�J6bP,`��c���Uu T�(�[)V ��e�^����&�9�Up���7
��&JJr�9���Mp;�=G����Uq�v��eR�e771��b����i��
[��W�߫�?��i�6<lh��"��߻���w��a����h�	M[a�� q`��L6�ɯ�T)�����$c��$�X��#�`rR	���n
���G��ϓ�{�j����������񝇊�o�k��~�tY�*�	t�h&/;;4;Oz	R�,J�Jk����*3]LM��[iC#��}�F���`�aќ�����l�-�;�r\�bY�mn���b�w�H�*�b��f���VE~�6�s��R3T����PA{q��䪤�.�6���ꋶ+��M*�A$�=� %��#T�r[1�>ة��A��������ڍW�%��b�Q5�ggζ��[GT��%���M���h��q	�]��;PZfX�b�J[G	aW�Ԗ�A���6K��u	T���^��K����HI��!9�Ւ	�2Ȱ8U�}��jzdԢ���*.��nu���:���b�Ǯ��s�H�sn���#A����1"��wG~�7[i�2��p�]\��q�����e��wQ�R"��<�.�Y7��i� &�Z=��cz�a�$�J�n��f4�jCb#�ʽ���J{<'?��ԙ�D��#��Cu@��
c���5�� 6L]}�
��ǹqQ���|Pp���O Z�d�z0�����Vv�dem�q�+�Z�v-)V'Q��\g!?}��L�Z�t���~ ֽ���y�H''÷�k>�,T
��B�Y�MIR�����x����gAzca �����h{ �k�mR�H�IL�>�>�03�NɃ@B$�Zr!u�|�oJ��ϲ�z���Z�O֪�ZQ���=������SW��EObi�0bin�DD���'�x�+~Xӻ���{�'	�M>��b��"�����r���o�.����� ����7�V-F��,l�1����}g�6i;/�!ˍ�B�7�#Q_Qђ9�Ŀ��bN�Q����P׽�^�vo5p^�� ����M�������@p�"�)�߮7�=UO��*/a,z#muRu�5ϝ>��?Sb���ls�<�W��g
�(!W>N�R������3�u$-l_�:�D�F�p|dļ�e�7 <��B`��C�7�և7�'�駝���c������N~�<n���T��)nv"*��q��`�p����1�� 
A�E�X�Fj�E/�;�X���>c�)�e�h�nfθ,�gH�-��@�UyVY��� �����z�njKݡ��� [����q�~M^^]�7��/�<�㒖��&����
X�A��
% �a�#"6Y�����|[����7r�gβ��V?��F���ǥ�5MG��/��7��%����'%���|�EE�����v�� ��x��S2�ps�O�&�n�����;Q+�ݪ����r�؂�z�\����)9�d�|�kd��[���o���M5�y��hZ(mU�{���"���Vod%����`t�E��'eH�J��v����G�h�E3y�$Z��i�N
b��n�.;��̟>���PU�k&�ل�	�+���c�}??�˗��?�t�1鍾"�mm�������;�P ������
ğ��j���(C�:����J	�0��$P�\��t����ԙXV�q��뫂l���t�̿�v�tm�<���u�ģ�/)�����l�C��d�s�؀Q�mhi	�,h[+"�}��ң='�[��-���u��#���K���dL����j|X����� o�
'�7ߑq�o���<���A��\�aaDS+Z��=n)W��������J�b���U]��fH������~Csj�_�Z�nɯ�̓�}�HFG��h�'�n��w�DZSg�̈́�I��3�s�D���D��Y�v_r-���ȍ_��@�F�xn|h2���f�)Ĕ�k���S�m�ҬFIR��2�Kj�	$�CL�Y,��M(Ɇ���q�Op>��QH$'%大�����������KH{�l�i�����dm���M�t����b�*�u`�o���(��N�L+�O��u�A9X�9�B�11�d�1ƞ�ᰬ�
9�� �B�0��қ����X�X9�������Ⴙ؏�ۻ��b#�&VVb'�8gS�Ft[�x̾a�H������Jg辱o3ԁZ�_��%^n���N 2��j0�}�G����Q��]�u�Ժ��X�?�?�>&iFAäG��[�B`*d�i�����DKγy	ʎ��.�2����(*�ԧ_��aa���%>��/٩�8}RL�HK$dBY�!Q�j�1�:o[G�X\o௬��k�{������_5[����xB�	���]�T�#uQ��7��
9Z����QRǲϒ!T�7��Q�&6�o@w���(�z_�����=�Y/k��U����h{&(�^�;qI)c��܀��_T�p*R���`�����3yu�BuW��CBy� �'�eO�>$$�1�:�]�C[��_^�t�~�6�O�*�rT�F����ńA���
���5̈��6�w���A�>��RD�(W'x����IxS�x�-J�HҾ��)C����)��닉�k{�T=&>7��`��N�)��O��9(�VW�>�>�O���7s�h��I�l-^D��=뉨�(�~:\_�z	2�����6`��oQ�>�����rH���tKȿċ+��&���ƍ>��=���[��S�W�@�7�et������wΊ�p���>a!�0 5Z~�޷�Y'�$��`J��K/�����}n�R��6.��q�<|гU&�d���� �f�Ρ�F	p&��j��e�*��t'�d��_[��嗻C��H��"̃3T�u;���i�M8�B,��:��ji@�qn��b-�bq4F�Gl�kD����&'5tR�й�?T����9P1���܎���	ed��V4(5�[8��U�s�t�&��Y5�������@3]���;��U�V��zw��@��!Q\Y���q�?��޹/(�
4�<Mn��:1��0�oϳ���Q؆�������M{�F	ѣ �����ɣ`[d��.�ڂ0�l	)��ި�s���ūu&������a���r�I$�q����'�h5~��&��¨.8>�Jc���a�'�oE2#j�����"#S�ܜ�4JW���y�a�j����2eU����1<.J�8q�]�~����YS������q3F��A(L'���:��Wb����kFt����=b~�#��C�%(VĻ���q��g�4^O!A��\(�}+�X� �c�m�-)�uY���l������t��g��9���'.S�b*����M2!��d�G=��x����)�[��� wj��=	T(sֆ��6�ͻ�2S��MS�~Kym�������5{|�hv�n����c��~el�kt���[���U2!JX����}�k\��B/�B;:�%fr����E����+E|��~}"��V89���yN�W�㢹q��p��i���Zf�O��J<㹤Iy�c ����t'/�7J�GQ������~�k�1���;�·�0�ww�JkIΉژ/��X�3��ߛi��F-͙!�>�����I�O�t�,"��i�2�?J&����y��.��_7
����Z��#*tǯ�n���d�+(.�>��W�ϱ�#��x����/x(5��e��N�L�؃Z�*��yTQF�^���+��d��c���t!?�؆!�����.��R��q3#c(�A�P}T���8�YÙ㭝}���u7�vw��X�OF֗D˯zRU]�J2�����	.�k�����7��d,܄��]B �7��q�4{<ݬ�X$>�9Ua�:�N�`N�K�Nx�_���&Į�f7nP.M��p���B����pJ��@���!M�� 	��9������d�h��`}p�xr�P�ռw����y��^�-D%q}����QRH�ӈ��z��C(�b�B/� �����p�r�=���g}f�M�{�9jp�R%'FW9h�@�DF>>��˽Pu������H���li��L�b3���*/�,=�{c'�ؽD-ë,"�cS]��^F�ֱ�|�+Ц��Ih2m�����y�����h���,�� �w^��(��r��B�fz�\�X��3�N�B^��dH�����!F��k��z�l�Ǆ��R�ﴌ��"��ja���U�_��}�Z0��͖0���Mc��˙^{o�j(��۵��А�GJ�6b��������*Q���E� &.��'u%���7���c؏�vv/�ɔ/�/�|�O��ws ��6갇x���՛�����d*�[��%�D�]u�]nnb�U���I���a���hz��D?���4�eܨ�YyɃ����OdˋriΪ ~��~�{��I�B4� �wE.�40�/����m���kܿ��S&Xw�F-��hKM�a<p��W"Ȧ^���"�}����1�ReT�B
�w��]h'>}������io�����"\�W���M��[�n�˅�l}��r�`�]��߹;�	,E��E�O<����\���Q�sC�ĺ"������_�l�fA�Un�qj��Uf��In�Q�� �U��WP0a��^�}<�p,s�V�	��QN�:��f1C�DV6̫W-����(+�,�������*��>s�W:ȉ���?\�I�� �j���NA�D��¼_���٨�-�TJ� 7w�L��jWey�Ue�D�g�d
~c�=M��8H�J`��o9����XF&Y�x�x'�he�㴾�;��"-��z����|R(}=JY�<O%�0�ׅ��m�V�� Z2Oy��^�ӸnZ����vQ�j���ǳ��=ߍ��p��?��r�t���ӝH��/::�7��6U�) �5�t0�fD4�p�{�N��h�P����Um���vV�0���}������])���5T��<.��XRL�wZ�l��^�ܻl�\<uu��hX�J@��aV&���9�ql���O�	\�:�vMM͚��@���䆸�t4xW��~5�{^��\Y�����X��l�LH�R�ꂡK�07_��$2��N�|��J��N�l0�t�Ib#��p�۵�o7��8Ml�y͟�b��z��VT�:�k!:q%��خr^��4q/�17�f����v�WB��#)&�ݡWj�/P|Ȫ�E�E�]��0���I������ʢ�0�_�h
<A����]�`�S��K!�V8uB?@^�����\Mڶy�m~^IHi��J
�����r�(�|fHt�5HR�,�	��Y'ʖ�$��ՓhS��9�ݹ�6��C�ψ��М�5���.��4#Z�L1��e�`�l5�r���C'��yB;�>׫�م*�s5~sH8N�b�W{�O(�ƿ��jD0����ݚ�c��׊e���t�k�������8��Q/�z��vRkk]�����7ߍ�/�&����Q�HY�x��J�g�Y
h���b��Y��s�5q_��7g� r��������(t5�|�@\/ �Y�o'�7e�s4h�'y�Fߛ��as]RXK����>o��B��k�"���2T�� ����/��t����P؎d��{IHx)�H��mYm�p��c���[ګ�sj���dnwP0�M���M
��<��¨�c���6�H���dm�Od�����kA.c�T�7o��x�p��E6N�Ş�)V�'x�E�p�����-����1l�a�t�.kS�ܦ���^�~�!��� d��L@�ߏm�c�R��^[�#����|�;֕�G˚Y�Ϗ��	�vP�GG��F�����O`���Ӕ�]�͓��NMO7����i-.�s��cǒ��^�@��{
!N����-)as��Ň� \ ���M�u����O0CF�)i�>_�Ul^ao�����Kl�*l�艤/�۶W����&�LT��O���n��Sx��YYw�{������7{�g�:\]��Qk�;L��=K!4�����5�[[����1�z�_��3K}S����Žá;��	�g��8Ǆ��_��/2�����ꨨ���CRJJ�")�-�(�݈t���3��"-!)� 9�    �� 9� C|g���~k}���z]�9{��y��y�~�9>�B�PE�/��~����B��z6=��[������YcAHZFPE+���m�3_���}/N��ɮ��G%FUY����͎Q̡��̈����GS
�7s�&Q�p�Є{�ڢ;p:�d�J����� ��U������>�V��ރ�eȢ����_fF`⧵����}�o�7&W�RF�s���8UJ"�e��yw�׳b�����i@�WL}�P�0���;��(2�8q"I�hR{��y��-t��P<m����BWUi���W$�����s_��-�}�<��jb�����Ź���\�h�OO
D�t���S�T���^S�W�eˁ��7jxnV�z�r������ؿ�m�k
%�=`�u@2���F~����aBʞ��7I�Nc���pP^�|F	����C�~���R[SWr|��3d�rN�.�J05�67w���R ��X����n���`����q���F���@�C��<�1Uk��?�|�ϓX1 ���M�7�=��k�\�o��>��r������M ��wk�0�����%��f=�pA_H#wO�p#����ވ�+k�(X�,O%%�p,��R_�c���׮vq�Q�Sc���*���x�x^��.�P%��41W�SE3���ƪ� �|V�|6�=��E&j$.����j�`a���z~�
��t��0l��))���x�Dk�T����k� M�ب�|{��<�	�%��J���&�~�H~u�{T�6�@F���u�c;Rgɮ�:i���Ղ���Ћ߼�pY��9o�o� ��Iɚn�UEg��Ǌ`�������f�����!I��T ��oë��bT0��b�Z�ݪ�}ӎ����s9�#klbB	w���d��y�'Qm�&)���/D훹�/���;*���k��w�0�����Վ\�.�k��.ڴ������ݥ*RB�<�@y�|`�����pa"�v��r��Y��������-X��I��z��m\�� �zgY9gJո#{�eE����*zi�G���:b����j�'!,i�p�K�8st)���.����H�-��E�� ?�9���r��x[ٺ���g>�l�k��t�u��O��l>�%|�W�j���lN�6�E�������i�i������K���c  ɞ��"�.�"{�Ȗ;�[���
����K8�/�����0ֶ��4j4<�M{;��)��# �Mb���~4�����`fe�nQZ�B�;�����:8�}^Q�[+b\.E��qN��k
��B����冣�\����-P��衽��r����B�:z.L�N����t���H�d���������#UN:>u����ą�=e]H����5�?7�p��Wa��`�r���R�Q�
;�x�L�SO��0BO��W�'�XXb��q~��#�~����`~Fێ�:m�.��T�*C�t
?��t6.�S��	���=��+#�q��F��`^�w��;�cj�s�;�`ȷj���֔��������oQ���o.椒��ZS���tL�9%u���_
�������<$�t&��)з ��yƯ�E��#7�j�0N#�sr�p��c�+����=*�Q��>��Rn�G���)�N��g�HY6S�Q��66lB��D�m�Kd&6)��'���YcaG\�~��A8�����9pu�5;��F.��j����w1�=L"��C���&cB��@��ZQ������-��$
"��y4��]�T`Y�����Zh��ځ�g�ô�LBɢ؄D��VY��r����y��w".�5x�1FUo�T|8�tLLrr|�zst`��1��SI��i���;��$^\^��� )R�C�%z��1U�&T&*�=�BW���6���k|T�l�Fn��
N�L�zg+��'�*ѝ���$<eB|�2�O����bK!�:Ĩ�WnOm=�����nɊ��5j�B~������v}ĈOt�vg�p�颫��iCa������0�3Ά���g	�џ��5~ĳ���7����t�"ID/M6��a$N�p�.��|��
Bl$���\1t$�L�!����	I�� b�{Z�>��ό�eX-�U��H���L����&8������	�<y����˅�S⻨����oڧ�t�� ����vt��#m}R���oB"�I�����{����JJc�ՁgV����|�O�%9m�q���8�k]f��Y"�
j>˰�ֲ�W$TV�*��^��)����I��b#��ސ�~�����Ol+���O���n~�L�74U���$�����ʫ���O�����|�*�[D��i�z��q�o�3���,c��#"O����/������vʖ+@�
bIket�������qZǙ���J��j8�j�-gF�Vl^(���ߗKJ)�t���]X؊�WJ, -��WѾwo�+��3s[lJL�z<>1n�1������gCw�tf�̆W�@����~I��t�_�nn��.辵� ���q�cĞ
�h�TQN��~�^4��x�}��S{�q��U����Q�U|ٱ��Wh��g}F�Zh�-����ܒv�Q��0�m|?�����g�Ʉ=9�͢��Nl���eˑ@�}����J;�~l�6qˋvdf� &4��J�+zä�S��ۻë��|���l��������u�$��%�����2����[����s��JDH�p�����Wǁ�ǧ�g2�)���% ����w�`*�5��j�*-����k����ӊ�?�lH��lU���ϐ����O�T�%����n}Ya�"a�#+�C�T�嫇�-`�،y��/�	g��X�1 "�,ʼPP����J����u�1�zd&u��]����95���Q�,�w��7/f��~'ݎ���b�a^���͒�.�>l^�n��Ȭ�fnO�E�z�A��2/<�	p���{EA蹌)Ɉ�c ɨ����O����k����/�*!�+XRĴ�'�NOFn�E=ÞbtC����ǘ���J�ts�5K�*�����CeR����XJEt(mgm��u}q�����Ug��
�;z�8N�9���{{Ka���>�ۺ��7|����d0D��HI�o�PM�N�M���]�L�o����Ѽ�nt�@{\I�'�Y�/�a��w�_E��Ȟ����_�B�5]�b���xf�h�;���Y��a���5ܴ�g��v5�'8���w�#��E-Y�	��WU�{��h�M���UQa��#5�F[����A�n�N���	F '����:����&�y��.\��0Hlr>�il^֮o�Wݒj��Lm�pf��n��A�U��d��שDad�2����Z�Jg��{ڣ���As0�;�zy�_���:�6���ɦ�5r|�B��#�<��$�m��&����K^�rYЌ�#�!y���f�Nɝ�tT�A\s�uּ�z	K����ȸ��ۉX�>�ӏLJ?�aS�P�j�&��^s�/��*�N��D6�w�v�]$��YŮ'G�����J�T^��)l�X�=2ʢ�u����*���VDm�	�{��gi���#+I�B���UE1���l�r�A���#w:['�ϼ�K�޾&��d������ϳ'������$��.{���/�}�9�C�S{�ZB�;g"�\�y��*����r1r�lC�@6��y�gX�����f�\)�q��ʹO�]%F�}|jW��1��ڒD�дZjY�`j���5����S�T}����ԀAU8�����?����΁3�=���w��W�j��sd)�7]��qT��b��HLJ�EE��}��I|�pÑ]'�b�_���.����PH�_�u{j׫"k}<��k8\})�'��U<p��������r�����(*��N�#�/�����th�*4n`���y	&,6��bVEa���$�u���w��N����ﯺT�2����w` a1"����������_ճ�,�=�t�1ޡr�=8��H�����t��Pj�N`�4�$��ǧү2�1�k���uS?cr�sw�ϫ�?�x��w��
"����~������z�Ycj��2/��)&2�'�
�'�L�Ʀ�����R�y��Z���3~��ձ��؈0�E[���8�֟���
����M��L�ݰ"s.�Ha�?̢�R/uNW�y�� ����Ͽd���t�n��6!�oRa�vR����\�Q�����9�n%�]w�Q�����M�Q�1m�
�1�-��5���ȿ�b�A���l_�F�ܵ���Q:u��n��o�Uc2�o�@Z�J�NB�����A�*��8���{8<�>��&�В�M��c��.?�B,g|߄�8,eN�}�X��X�?j������Ak~�o��a��"�X�{ ���`�������з���K_a�B��Rj�����f�yO$��; 
)VJy�C1�n��u���Rs� � ��ox���sb�u��E�b���ZC�O��N�{���22�)��,����(�~f��{Bʨ�M]6/Ɗ/�H쫐1��=�'K,��=���tv�q^���r�\, (�gIs�Ѩ�zF�eE���(B�ʖoV��P��HP��\w���-�r�6!�;8%���\Yg�g5:;���*��QD�$Dd ��@�,��l��[!����EIgf��ԝږMޝa,�0�/�в`V⊪ǽ��4�Yسb�z�+O�F��q���J�c�S.W�6���ΟL(�v��{ojwS�&m���F}{a���O�Ur$Ȟ�����E���1������%yr��1�����N�bN8�W^L$o�ǘT�����	�G�c�^Y��!!H3�Ca� �qz�|�W��o�+�;�U�:���w� l����͠{�����
 q�N{�q:����t�k��cf
"D依Ea��VU��z�	\ȑ�h1��1�ۻ�pnCja�_1�囱gO�G�L�<T���0q2�+�/9�V���$�$3�χ[]�7/y_�:F�FF�c�}d!/���z��r3}��vGg��z�ZA;r�Ǻ����[W�K5+^��zPT;鸬k��0������j��Y��l�c||�ar�:a�r����� VW���zaj��U2�̱
�=��|Ӭȼ�hb"�@�^�Fm�0��"��!��QR�bE�Mof�� ��l�5orB�W���6����I;�G�����zДx��
�{p�M���Xr��
�"u1C�]|Z��|9A�2�v���`�)1�-P.���	g�%K����g:X�ь�>,TU-˔������M�4[̭*�*,@2����ah�U�qؕc���ی�7&z�KiK��M<��8ڞE�t�=5H�E�|��d�0��y�-�W��s��{�6!�|��ˣ��� �p$����1 f�✦ �@J���J�����;*w�t�0T�=�wB�_�wڤ�I��7�R�z|>���� ǹ/���|�}�E�'t&5���l׏�������^^�x͇u�+l��U�y811��}�r
=��1���w�t-0TG<�7�9Ѓ���ic�`���>���S��`ⱖ$���u�Ԫ�0�xo��M��M*����^p�KH��;���{�L?�*���&q���h_)�V@�bǏ�2e�۸lc��K�Լk�[>[�>;m����9i0�r<j�K{U�6ѻ���bγ5�5�G�l5���ܤ��$� ��vh]��d��/��둪�� ��RXׇ읈��.��s�7�[��?��
M�ȍ���g��Aw�u�#�4�~g��Tk����>E�Ct�g�8G;�����c��x);�ɘ�������x��xV2Q�9�$u>(:��
��U� Y�NT�t~�r���F����@����H�@�^�_:���n9�;����L������ڈ�_��4�!o���KQ��|��しoUf!o�S����ӺeG�n����ӯH���t�����R;��QD�}��|��ba����/��#amȧ~�6�f���ӓq1ku��M��/�<MJ���:�.�Z��\s���͉��e�bַ���v�����H�g��n��ϲ��υk3J��#��`?������pw��.{XeTe1�zz�R��̢�@P�Jg��z�իN�\�b2Z��,�8�1_l�^�ϛ���wRBe�d�%��ѷRR�L���Ժ~�čǘ��x��kG��Q
�����+� ���8ʐ?/�M=)g���,<��@�Y��B��������r���ݶ�B&�Ю��WY��5ϳ�k�@-Կ�� r�N��bd�UN�Օ�c9e��>�U�S�M�G*�I�Ŏ����P/��k�䰟~8'$�:1��wRΫ���\\|���#�NkLo��������?;Sܬ�I)\ّ��Y����n��%����}�庡`
Z����S/��Qi��F_�z!�-�<�A˴wI�����s�S������l�6j�s����>��p&&
J3�W:M�$u�2�k-�cn�bO` �,���Sz�3�;�W-_�\�'6�i� ���x�s�F#�1�e3��:���y�s\1&M�`�Z�w|�n���m|{��ԗ�����P1O��N3��3�GR�Ľ���@�����1����ˏ���� <��AI�\m���b�}�K.�b�T�S��g���(;b�~~��>�;�����F��߶�����ep�MH����<j�l+5EI��{w�i�A�e���Qz���,�|(2_�0q��ycڌ'E[���+�U������{~��V_�u~L��(�]�+�����w�d����%���q'm��`�+^!q\���Գ�+��%*� ��Ə��/�N�Ο��i�=@gG9Gu� ��p]�5(�Z��Uߟ��©��é9�M��&i��g��3Ry/��w�f�v���[u�������A
����>	�]��+��g�|t#G�Tk�2�p��NQ5�_{��r8�H���=eװ��NՁ�23��q
�J���K�/�\=T[�!���T���tA��S6�bK$gr������J�y�b��F��k]�gj�
�o�d�#��HCcq�>��U��Ԑ�M��	
�������x��-m�|���^���kz�A�k�t��d���b
Bk��*������g���2~L%L��\����j����$�����H��!A�T�m�ϡ\[�z$L��J���\Tz�:Rc�����LƳ�+�lK�J ���3z�R(�>�,i�+\�SF��o�yD�\���=IZ�M)A�"V4�`~d�e=�Q�ŗ).�%������T_��Z�~�Z��d��"2�J��N�L�ю(��k����S� rașTy��R��z�l����Y*2AJd���tZ�(<[䓰G�i%�����N�N3�-p������]�@fD��l�ʣO|��v���� ܇����v�d��6����� �k��)���"��ba	�3�gr�Qҥ���1+���7�'�1z"YT$˾^
�ޗ�C��ֈ�77�%n;'���LHX�0�5����փ�#\��?2F��Ea�`�E<EE��8'���g�t���������|j�UCra�6�kNV���.S;/�#��'�������:���;�L����s�^h�b��ՕX���G����eϳ++�]Q�A��4@��	�:�ʟ)o���|H"�>m��A�I���,�^˖�[/���j8
�T"���/�|�$��͹��2ڏ�Y��Z?�;e��Qg��4�nT0�_%���w� Ỹ��u�Nc�%�^�r&Ϲ���i�|+�n^�G�)�&��b6�gԌ���Կ�7������9X~Ƌ�1�3ry�Mm��m��K��8O.�#�;n�4�tȇ]�:3.Nmߞ+x���� x�<��v&<�:����v�z�߁ؖk	��9�^]7�l�J\O;m��3�t7�;���vw�4�ţw�g[��7p�+���^�
<Co7ST�lix���$0Ya�(�F��X�D,<�S_��Uf�vA��i�B3�Po��H�/Z�����ŕ��-w��	,`��ԋ�J>.yfO3O�Y;y�zI��[0}گ�GU���^�80i*��[>*�/���+\� ����1P�l���ӥ������i��p���"ے6�П.����L�5]�t�� �6�<$n�)m�/c��)���G_���X�ߏ�w�:�=�m�d�'�.���������着D"��)h�<"�%���N��hh�Kq\.�ё��o�(�Z����䋞��mww�I�p��xֿw$`b'ӛ�6�o����4��t�Cb_5�j�F���N8A%=�h_p���5��-[V!��-Al3�ٍ+)��߆�gk�Qawvs�Bg~��'m��Mt������}�>�1�[0Zb@:00޸��p��d��ϲe� ������k?a9S��/��e&�����.>�)"�B�h{U�`e���k ��V��kk!��-�� M�Љ�cr �>%�z���o��j�����u��,��x��ͥ
�4J���n}v�v6/�ʎOw��,�u&� ��T�rd�;�	1�-������>��o$(��y�Vڨ@ޓϲ?����F��w\	r�{ LgMv0^��o5@ެ�\�����!*R��9�g�	��?LM	_3#�ƑKǧ#b�mz��y��ʀb�o�p�	=*�@����5/�c���ۓͥlS�	3�K.�7XS�ү�9���tTAhu,��lNԟR������n�;=Z���ÿ����R?��۫D�@�?bm� 966bB���aP���)E��_�!��f?[�X��{�S��e�u=7kB\��*�H�_%6�M����0���eS*�C@4�J�R����Q��B�1�9a��x ��i�
�ߡ�} MQ65E ���h��/��a��;����{�^"����΋�/㍅s��e9$	A�&�AM�UU����-|*<ch/��T~��K-����BoPT;D3'��O/vbq!��F�����M�BN/��Oo�O5��BG39v^Z<���������{<0��Lb �S���D�2��4NP�R��F�!$�j6%���R����<D�a����)5�Haӧ���?pvsT�M1�ФF=1U��B�5����ݣ����3(��HU��p
S�l�(�;o㎫�|�-�N��(��.����smT�NN����YK$[H�o>�m$��4A�C@+$��r��ﷀ80��44t$�wS&�����M7���Sl͔�k@��'�[�*O��0����6�G$D}�B���Ћ�^�����Ɲp�D�����4��$2z�W&��ZK����iX�G2<����%�!��m��@f�4����Ab�q?��6^��ז6 W��Hm�d�B�}�W{,�U�  W
�)�ץ��F���	�)H����C���DN�)���g~�
�n�r������K�zğ{V(�E�J+��[S$�;>�2ܤV�!��|�n�ǯu�20`��йR%�7O�J�<��vT������iEʷ[����gk�{
��<�{~�Ϯ�;�n���_]}��ߝ`L�W!ߧ����x� �L��yT��x�����w��n`�d]�U�r.���)k�tv��n��c�2ڏV� ��?�"5�6��:hŵ���q!��ԛQpp��
��[c�V9��G��cO���ߏ�ʎ0��[�ޫ�c}R�ȫ��Y_� F ���Ϫ���NA^�Թ��`�BtXA^�B�h����B��%����y�J�=��)쒱�r��"�[�9��1xt�r�wJ<�й��h�:���iW�p�9���YU�A����t��ªc�����?����p�Y�w���S�e��i��t���3�>�q��f�-8/q�����S�zl�.��"7�jEF��K��#��+��}�>ݜ9��t�6R�J�ݷ{�����Rqg�'w���@K�{.�@h��sr^�`aBf�&N~+(�[����P�����c�\��{12�H
��@�j7�������i_RO�)�̆y�=
��)��Y`��[{sO�(�O�X�%#F�6��آڟ.C@B��
��cMZ
��#3s|P���	8M���VXOʐ��^�;\�Ь�$�8�ͷ�"uʮh���z�>5�/��ه\~�e~_�q_����z���?��<PDۈ-��EvR'���\8}@���,n�_X���ߪ7`���m��v��/���n�ߴ�d)u�_�EU_D�����Y=��ˑ�X�c�u�}s��H�t<72�p��V�X�u���p9����9hu���� �M&�p|iȝ)o���`�Zտ�DR��`��Z8́v	�mkj+=r�q0�Y�<P��h��Ňp�m	��d,Q'�[SΈ�s�"��}I�����%�d����D��S�>�.F!ї�����'�\���@��p�̥�&A�GV�kkA�Ʒ�o����&$�I�H5^oo�ET��K4��q�7�nKmѓ-�n�p��8X9�k6��yi��h7w��?�i�ЙKy���Kr	��[Q�-��m�_�B��Fz}#������� ۫���A������ܕ��>�_RJhb�iȏ������VP{6J�+0/�__�O��f��Y������&���"��cw��I�>o��HШ�ۋ���Eɕ��H�j)��6*哤&ѵ�`/��1���):�y�yW�p9�����e6�z��GM��y��S�ͨ���,J�(7���[���ۿ�-�iͺ��V�BrU�G�VΝz ʴ�w+y�CZ}ՏQ�W��+��O�ߌ����CPQ1���D�3�aX�ۤΌ�Y���زd;ܠ$�(%
�92&n�e �OHv�tNT����r��h͐�ԓ��x�`_��P�Ḕ�1����*����` A�)>[z�#�g�#c	��^-+Z jd�,�� j5���L�H=A��]�'k@l[���a� roW�����н���i4"��Ƽ�g0.�w�&r��) �E#%��69o2��u�画0��-H4!}Ɯ[��L`��/���[p�ap�,�L�lX��b8#c����ZV�I��x��Q��Ol��Hl-�%$�_`�}���ܬ�X�y������硔ܾ��~W���c����'5��ӭXV��}���$�^��~��>�-$�=I�2.�Oy�^$ KE:OF��'ٵc �5��2�@܉ޏ�Ы�fm;�����T�mH$u�S�y�ү�S�|�Q!|-^�`Cb@.�O�~օQ�΅��\n�ն�!��� ~ H�����G_Z�/�,�^��M�3���#�g:S�WЋ�#�#gp���1)2��������`�Y�L!�����;��ͮv�ՙѮ��4���!�cD��Cy�h��/�E�a�L��b 9H�c!��=���n���e�юq��l)��5���������􏩃Ǻ���b3�@_���?i�������Z�xR�����R�w�>�c"���(�U.��푒&��.ZA�1qD��;
h-8�V�$�6!;�f��O[-�<-:�ͫ��\�g�ƒ�a�<]7	&X:����^<��{����{tBfq�eM0Ú땄f&*�TW�u�?� ��R��8�F���mL[�67t=�n��cN�����D����� �-yQ"8w+�y ��H7��^GN/�@&��emS�	r���J��mU��x�o������ ��o�s�W���	���qaP�c�� -Fn2��ꍚR;����ށޔ<j�W�4OL�HLZ
�������b�j�b�ni~ΰ�3���2�\l��l���[�J���۪C����H];�;��  ���AWװvWڗ����%�]|�3�����^�][T�v��7���_j�Q'�g.�3p����9��v ��;5��'����oIo���ؔ@�14��ǿ;B��i-O��ׯ����X���3��z�Й����]��p������$��3�^�{"|����j�[i�3?g��;���o*��"�م����U%%R������6�nc`x����IÌH�ו﷈wHpo%�O�@��Ҕ�� D�;V�.d�C�%��� ���dŗ���Q���f��7�<�6���ʣ��-�5��]P�jgD�K(�7�r*ͥ���z�}��zc�׌�����R����p�x�!AD�=���Y��r�Z�ٶ� ��г���"�32ğ���Y�j����)#� ����'��ک�#�G�x���~�!��]Q>�7L���̣J�`����:*�'��OM���-��çV�.8�#Y�Kϟ��[��_'m0�V&`���?j�,����ro�f3t�]��?dz�o�aO���Y�V±r��h�	�;�1p9�֜��%��&�()�e��?����.��j�+�"D����X���P�8|A�0%娆 ��#c5��%W�v�%���&gZ�+�H�q�� �e�[5��%I!������P>2gĜ-d6��1��C�;K�JsK4:��Oho_x�m����q��afv�#X�O�ٟ��m���U��)�I����Q�/��`o^e��y����5�\�������; �������P�E���Ku�ׂ�nхsa�t����0�ސJ>5f���.n�N�֐$ :��셈�*\��x���L8�Z`Ϛׇ��9��2ľ[{��<܇��2��07�:%��T��Y�G�fR��.��ES\���B�Qh툉��EI�痧���»���m!r0���R��iu�ϛ��q�@7�pd�q�ФQ@`&�j
!|��*j������Ǯ�����u�V����r̲<<��Hۚ8�O`��{t�#�85��/��ǉ�8��A����=_���1/׳pj�:O�� |s��o�d�.�^���77��&+Z���SJ�ƴ���J���N�W�R��z����''�O�X��P'A���n�۩�Z7��<^a��I���lU�����k:���*��Ȟ����P��=����Nj��GZ�A��cՀH8�=ݍ�QBb�Ao��L��cp�X��EY�.��=Ø�g>��O8���L��l�`�	���${BW�����Kw}D�kZ��<+]�Nυ���;]!["�Ϡ��B@��:�|聘xE���+)NA�r(�s�=58��1-[!�Ng���1 H�'��|)�M�����?�b����YSN�����1�vEx�sP.��sPZ��x������ssm�l����`������xr�o-8�<l�ɦ�}{W��LX�X�l,(9突:�o�6����#��kF�R�����q��"�r��2��	�h)!5�!�" Of�&y�� ���\���V����kd^z��h������A�OK&�B�x�k�A�%)���C�N:[���A�1}H)MG���z��X#K(<o�c�����ж������0qՉB�?�[^����@rYT��Gc)u�-3_η[%�F$=�����s7߹��զ�]��n���q�:�u��E&X��|ď�k��*��B��>8#[ջ�1&$$�;6�"�.a	���
2���kO��ft"��fe�~4MS�S{9j��;�����bn�J�M`9����r�}��#�+i.]�����>��KJ%4�ZJ�?C�1���QT��@��>�l3�~��!XO�o`
r���������Q������|d�2�x�����(�6��V��n?���
y9�F��"g����΁-x�q'�B�}��烳��C��HA�������F�z VAΥ[�4�#)�����at��@YT���������c����f�G��vD�b�����xI�`�[�4�i|��x�{�;����U������kC�Ho��FNj�������6@*�"y\��U�;��4��Z����i�g�N�oJ4	H5�"m�,MG/��^����^����v8��~4�s�tL\^ϔE@O=./p ��67����=���p!Gߞ�ҹ�z�N��Np�i�R�5��)�5���#�fC����uǅ4��ʈ;y��]��s�0\�n�܅Dbp�u
a����Op�9c�P�����@����p���⁹�K�Ƭ'NꍷF�����V��,i���X��`\��rj�;3�W]vU��*? ^=�����T�����F"�ޒv�z_����DrX?�>V�����5o���~�&p�����Aߺ�'R��p�"gL��gB�.o(��_i�<bM���F���B����]�]Ӯ���o�X1᫸�LD�V�+������R�__�wq�U]�I�2BB)+�{R�<�Μ��]�x]�H�nBm]�����{�ɮr�h����X��H��ľgƀ��<��,Ϛ���R!��+X��Y�d�9|eG���s�K>!ê��8
N�k��-�� Ζ�󭬞�����Q��1g	.�R�l�*��Z�U»��� ��a�&Xv_Y
���|��&Vĩ0O�Bg��Gf����GD�像�Boj8��8単4�J�͋��L��)����3�=��,Kd���=����_�m�Ʉ������H�_�"��:�p�y������c��{Gk:tՊ_ޞ�"�#��)����M�{V~HZ��׋X�Az,Hl��1c�߱���If�G�3C�t.Ժ�U$�7���͖(��ԈI���8��$��8f��ԗ��_�(��|~����e�OG�Eo$�e�A�̼�hs�&0f��pF\\k gq��t+	��J������0+wA��@�]��h�s/F��0a�8�2�R�-j�e�X����x�ѽ�	TnՐ��z��D���w.��rR��L-����@�ĳA�͆����o��]E�Y)��1��".�t%���c��4�b��0����4��8��"�rpvt$��'%��`������_�:��#�J��V.�nY�������N�q�?��L�7�P-I�`B`�N�:~l�,�F伡.����#�͠ �Ws�|``5幰�])��f��Ø���t�&u`�4S ���U�����}6�7��Ō����*�G���Ƿ�rᓭ)~V�'3 �"�F�0����Չ���@
70���~ȞJZ���j�${f/2V�xﲨX��j~d~��_�5ԭ��΃�@�;�^�#��|��bs����/�����B_r����;.h��v�����7�\��T�$Y��I�Ĳk�[����D;����2�N��ͳ� �u�՘gAg?R��t�̲?�/H����_}-�U郎�\���S���*��.�w�K�հ��쨣�ѷY� ���Nɱ��4}�b���~i-/�d�^�Qͣ�(uv��39E� �����5�6`�y�\���P���+�i����??	'�IP�M�����涚�eּ��,P��ޫ���?c����;�T������z�v� ����D�pך���x˙sy����mb��O�<��i��>j�	&�y�^�N�بgk���$�t��7r��J���\��\�յ��KK�
M�{33MPT�<>^���@�ۯp� ����%�vf[�)偝Ebb��o�ž�Vb��̏��W�\}�B&�'+�Bx�a���Ow�Ծ��o,�������M����G4���
ڝ�������_0G�����"��<�Q�w}g�Py��?�ž�h�sM�z� )\��<!l��B�װl>�z��PJ;\*r�ߋRk:?�����3��	Zm
{�7�1?����̱ٙ�ة�LtM��[?I�/h�W�jI���@�u�;�5Ew�z
�^�� ��S.}%M�6�)9�w��}��$����o΍F���LW�� �L�zń^z���P�q�⺵ԕ�+H�Ry���@�[>��Gv�L[�(�g��;q����?R�G
X�-zE!^>�K�������{�k�q����%e�1�4�Q��h�k�;��A�:�pb��l�8�8dH+UM�O{���8(��sb�G;b�N]�o�l���>�?]�[���]�I�(��Em ��i��G�\���uc#����U�F}�����b�i�Q�>	H҈ɅA����
*�O.<|�f����������8WZ����2s�^��ptzt��xؒ��/'cY��z�$���x��\�����嶐�G=u�A��)�����A���oȵ��5����]�7�
�.a!��X�N�I�{��t?�K�;;x�hg7}��2ᐺǸ��ׯ&�]�oG�Q7�v]�ŴG�%�U�i�{Vjp������xD��u�ErvR�Y�� `?AHid�,�� R�~�I]5� wEu)����^�u^I��V���RHFM��r�R_j_�-jyOW��U�k��W��+��5�=���X�l@����ۏ�1�J�C�o������a��l��d���l`�B�{-V+;�
��L��5��C�3愴����Q�W" L5EŽݘ��U��w�/�%�4_Y1��s%7ކ�R���0�I��^V�L�Cu{*�v� �g�+��w����3� !�� �c�n�r��
e�ـ]m��m�Kx�ir��Ŀ����%��`�#�@,�G�!��tEvYd�p'_2yh8�q�q�����HA�P�����tF]@zgΦ���g��&,��ס������2�i�t�L������mt���x��$n"CsO�e��!x��CWdU���C�Ψu+���u��%.��8�7m�i�4ҿ�g��<�)����l�o$�����K��a ]�����P��t�X��2��q���*S+��]���m7����S�&�'��8^��Q/��x�1<,S<�>T�5�^>�&J�k|̻�ru2����m<�2{�ǃ����mR�-���Gq�{ܼ�������z�޽�%4=[�[98�h��W4�����'����f���U�.O�%�6�4�56tL�}�n%� �̶����m�%2��筰3�uX=�$����k��iJ��H��ۏ����V�z������:�3)y���$^9��g�x���Q �3�;�3�#F��΍�f�4^�;5G��;k9%&�> y�#�h\����B��W�}N=tx��
ĩ�Dj���
qa��&���D�����aM�]�p\��Ea]�""J�^�G���ґ�Kh��(u�5�D@@@zOP�K�:��BK��L�}�x��}?���t23gN��}��Mfr��2�Tl��zΉ}^�S�j6�u2alr�2�X˕#��������L���'�t�@�n�ʀ���iq���@>Z9N@�3���6��h?'�Ӯ&a��H�O	����a|gO��\E����ʇ�q8X�9���*�R������ӐC�1ev�)����4�X�o�9�K	���!
+�WoO�l~"|:?p�s��Y�ȫJ�{�4��yz2+��^WA�
eQg���K�wE�V�Q7����sH�._-'��/ �^\�5�󹾯r��v�yN�>{��M����Ҍ1?Y��X��"2}[�~�ҭ=��t��f�D`a���՜��l.��-s\QY$�KJF�٢�ܲ7j�Y�����8���*��]��zz�.�yM����=����tqV�����v-���x�{6Z��ʗ�̝V}�A:�OfV��>yf�c��5Bz]jm:��ܹ��|k�Z㽫�n�� $>}"u����m�����pFf&�;6p�����Ȍ�{%�2�&8��!���a>������R�c�Jv6Jv�dg��Hֵ��d����3[U�`(�gȔ�����������fz�� Y�E���N<CS����=0���s��~���q��ʵ��Y?\i�u�w�*�8`溯8��`�K�M��ޭqT��᪡/�u&]l_A�X���e|Y_=i2Ns��i�������Hc<�n�t]��K�Z�3��9�;6��ǳ�'>��:χ�,+��ȶ0�~"2�8��:.��R-�2�Z�#��|��ҋ���+�o��6��l�>/�Ђ�w��,��}�A�@�!�xb���c0+$��:�8�Y���~����1�=-�V	���w����%u Yx{M<�2�j%W}�{:�1���d9��$ĕ�X#��²��:+��I���B�</8��Ռ����ȸ���y� r�O1��d��؜�L���fzg�~W��,݁>&�~z���#^�5G֐�[���#6{7]^N� ���w�Vp3�X��Tr�Oʫ����z�Z#95kē
0�镃�	?�78P�==��W��3us7�I�ە�Z��?qM�"_��H�O�e{�0f�t�bf�`f�����pn�����/E��?�e��z�I�f���wŗ�@:��N�r�H#�2�TJG�|X��R�O��!��@l�h8`�BL��e�vC��Yi�/޺y*n��)t-��₨G@�1�1r�������~�ͣ�1��n[��Vz��T&7 M�o�2fr2f��4O?��҃<��*k�j�D�Ʒ�_)�?�E����B�?m����z�x�TNn��i�N+p��%��m��X�>��B��`oq��T��l��F�nL�6��N�ʗ{�Én���_WۡBPg�����6i堾e�s��#e�Yj������E|�*m���4G��ϫ-��;�$�;p¯[����ٗT%���c�%��P"�"cNwbp��K�����(���E=��]8O\�������������嶟��K��b���.�7�����n�j޽k��Ok����������S��oz��jߛ6x��X@?���t��E9b�3��Ҏ�������S����� 4�}�]�7��B��A��6+�&�О�[��] 4��；��c�T���ESx�
��
{����Ș�Y�l�3�Uos���w:�^@";S�k�q�쾮@�X^dK�OAt�����]7�(Μ:����C
B��ʧM���)�a�����Y� ��
b�5�j�8�	�	�SW��C���� ��Z��^�b���•�L˽��S�N��'/ĝ8s{j�	�25z�O� ��3VR�������G���@J��:ޯ/g0Z�'�4��*܍)�`�EY�`��?3��-'�k7N�66�)�z�uQqϯ��"���2���ϳ.�}�d��e**EV��	� ��t* C�W�$a7R_<�#!Z��w��l\]I�g�	a����o�@J�X�vXLt��R~����n-k�_?w��K5X�_����c��>dx!�R/�qt���%��ޢ9crc��r��������ڧ�/Zj��|��"U�g����"�m�%Wֶ?�nw���x�v_��.@T��J�?�ܟC��:����3�ţ�|�Ej�F��#d[�孏�|N1���,�v���gw�l��!�<ǀA�[�=�9m3��Q;ϙ�G�f���u���A�|m���;=wý����3`�5��`#�qO6���_r7��}()��cOm'��NO|���?���U�滥fvZ��%�1���� �Al@�  J�����t�5o��V� �˕6p:���Ѽ���!��O!V]�jN9m�� 4m5S�FE���J�/�*���̖����n?���Q.��kk̛�~ԝ�H�Z�����b_N2�^엻�"#)Ȟ��p�˷��F��>�x��	�ష����u���R�(6O?��7��+�����L��Ypv��*/gcO�O�kU'�UY�����U���2ڂG�����K
�S�b��r ~��Y��u\l�~A(5]�퐡�[]n}Z�qʒ?��
i��`RN������_��i���,��yO��.�����=Y'��9ؕ53�n+sU�^�;��p2(���Ĺ��8�q�sF@����'W�d7;�#dw;U�r��i�Ͻ�erxa>$���9@���yOy>���ߡ�݆S��h^�hx@U����dV�R��H僘V}�t���ⱖ�8Ks���E^��Ԕ,r�7�0���|�W����2��F�������|8o��*��덻"�F���I�Ĺ�P�l�,/��:��S܈z	�̒t�×���\����9�d�5z����Լ;�q3��sť ۵�����8���ŝe��D6,�������|�Pw[��T��o56���khRGr�H4�m>`nJ��G)��`����:�M�;М/lʏ(�RQʻv�@{}�4Gs�9P菇�2:�I�ͨl	㙯G(��4����z��J�j��7X��{h(gF�[C?��8���������Y���![a�%sU�Y*���ʷZvf�oL�c���m����%6]��Ļ�d_ҟ1A����l�x��
'�p��V�KŴI҂#�-�u=���'��f��R�͜�]��6�2��.�;���w��
hFH���5�2����g<}���~x��#v��t[�K���~gR~�U�}/��/>+�}W�4�Y�u�y���5��*�@?�3��P�ZcՙW�`� v#@dn٦����ZԢ���.2�:yq4D�c���2Ax����Q��7P�ag=�Χyu~.�7�a�Q��Ө�]x{S��M�۩� 1�q�+ot?�Y��c��t'-�#������k�]S��
�ͶȬ�N��Mv��s��t�n��R��p<\@^\P��
��������a��������Vk�&��ai�]�H�5���[�f����L�$�� �xb��;���B6? C�r���L�~�hG
�"PZ�<���fo�Q��2�c8�2��D�)��X�����=I��vo^����S(K�[Ăm;09�M�Tr�<*�*�T{�� �|f���&��j^_w�|HY�c�j��Z�l"$t�D���j|@��~� ���'=��r4�b�.A�!��#x��1縦�\3.�#�R"]�����?(g`F�l�w�k��+e�c���olb2�B2	��"�שB��g���B�����$�Yce��|@������,)�\��G�w�zw�X�T��8����'¾8�H�}ac��o���cL^�)��F���|檝Y��r��G�V���ņ�[W-W]kO�.u��:y|<K-7���ty�Tw����`ݟV'ơ2<v=�w��PX��������(�^��q�ޚ�Y�����lRl>s:����Hb�g]3�bsn ��p#��f\zO�N�O�eo�0SH����;H.� �z �ƎeS�E1s"��2�~��e,qi���̞7z�����9/�����W���<,b��4g�	���R��Y7������3~�ц�h?Z�%��b|�m���$�� �����B�d���Dws��ak)�p[1�Mz|�J�Xi��=F\Z��^�.�!.͇��(��gԷ7������̾+8/^�k�q�(����]�U�TZ�S�l���PK����mȼ�$h�'�g����=�`��q*^����N��d����	}�;!���A�U�8ǘ6ǰ�:SY�W�=cf�{�]8i����@ePl*&ȇ��n`�J.vC
2�m0��(�hbcc;����2�?v�%J�i�'Ԏ����Vz��x�3VVl��f��Jn;�[��w�5BQQ���Ѹ�:�t,�~Oz��}
��͘����̀}�sY@�4�Q���$ �ݣ���-�!�1��i�J0bR�^�Ɩu�!u� ��=,s yI��49�"(Ή�ZtU�뫦��"�k�������� İ�A�W���D��_���mݜ0�z�{�9�G���� ������j��gj2�����l�j(�۵��� �P����̹[�܇F[W�.ܻ
��{-]�� .��MO&2D>�5��Z_-��>ӂ�vE���	/��|��"堬�Ƈ�v3��F)E��Q�L���F� dkvr��1A_�) �������'����X��@��p��'Ov���;/�1At=�-U,tk�� p��+��.l���`�"�2Z2֥�h��$�Ǿ%�����=���=�~y�?�̙��������%Ģ��@S���ӛ���>�J̚Ԛ�{f :Y������+�DiP���W���?���AAt���̲��4�C~��C�"�湛���ư����[͉�3�t�_-����ô��~��H�_�$��l�h���20K�A�&n nV%S�{��}6�t����SPTf��<���Z��I����@t�G�H�y��DC�GȬq�jď8���*t��D3�/gfg�i%�n�,��ک�w3G%�n���|([�f���^��9K6�[)����&�F!���\�N���V~x]cq%"3� �ڦ+�H�Ո�x�:#w���B��E,�,PW`��R�����^�᭍�l�X`��S[��'0>=�����f�I�����RĆ���u_Azgٞ��$����{i�[s�7{��17?�|��"����wF�!�������8���
M�W����:So�7Dǫ_�M�&<���eC�˳��lp���X��S~������Ia
�404��|7�1�KXR��TDD����0&�"��(/�X�qQ�Wm��u�!�0�;��
�2	�h8�\�� �lm��0�ww�S08�1XL=�a}U�;�S�뇭��9+���K��+��F^�����˗�{=�:�Lj�
����oЎ��N��z�����$ō�j�;�Vi\�qJdF��"�[����
�� {���EԚ|�[�ž[�	Ӿ.�G��n��KKp��,	~% t]�Ҹ}9i��L��b$��b���m�2|�@fв�v���5ZfJ�}����T�X���u���B.�fl��5�c�3�=\êӃ$!�Ǽ:
�;��T2z�W�~��RZ���{Q���C+��HhUV�jʲ�݄h�s��׋L��W���bh}FC�V2]�I��&�؋�nĨ�o�qpP�Ɋv��%��b��P�mu��Oܙp)�IrKr��SFG�q�[>���t��������0 ��9�����e�J��[�4^�\��0�c.�Q)�hoʥ�?661t����
"���4W���?��3�z�Cxnжp��܍��Q-��_u]����4s��w���10�v��՝<����@y�e�#LW�QgΪ�u����z�J5 )�g�޹���g�*S���I>�Q�N��C_z�3t�5��8}�|f��ጧTVM��=H� [�R�\w�g��_���Bޔ���G=_ג8�E�RZ�@0~�W���&�����~��d�I"<�su��_(sų�Ӿ��w��K��`�b�H$[�N�l*T��f9�͚=K{����
:ss�5�|��8K�r9#:�Z�����y_H�H���Տ��z��6�W��QJ��/`�Aν3F�B6/��� Wj��u�'��t��
���� r�S��MB�+�J������MJ�R��d� ؓȸ�\;{V-B$L�ӳW;?�EQ1s����	~�<Qq2�lrs�����3��3�[���q�,
(�����2Kog�����e�-�ǹ���k������u����;`�ǻ[�(5�c
���D�C���]ͣ$&��
k�8�v��3�u�ϰZ;h_������t{��W��	��H��Sb��q�ga0z?^��A�s8�w�03�ڎ2���ہ1�T�*���*kP��P�
�z�48��.ј���t��*aO��[��H��-�9X4����;aЭ���,�:*�,����T�>��bY�У�GYl�����&�%�ǰ����{c��XU�ږv�9;�9���ip!.�')�֛��s]c7����8g�QU��{7㙆.i�
4q.�P�4JBWV��| S��l����Ϥ�`\��M&�n���i��%MW�7�������>�3{#<��\]�c��M�@�/z}�OҢeg��A�1z�,6�57�V?��C����q�?6��6L�+��N�'VGA�oWj!��Z*HP��S	�$b�2��o|��s�DV=f�9 wBe���8� ��ۜ�í�4&%���~������y���#�>@qډ��Πǲ@XfU�u�ស����YOAR�'å.�11�>��L���0��H�q��U�C'h/���AN��OSO��������dxM����(!�q�I3���2�F����}��=54�[y���{�j�z��C(T���B��~����w��Wed�Ӫ���e"(YA
r�U�]@���xV����6�E��i݂�P���P��B�"�@��Gg`���� .hR��� �a��{�n�|�߂�z�ޑ����◲�;��l]0�=�T(8O���$�u|��J�� .�B��,�[����W*�
�}/ۘVPQ�fmf�8��(b�=�=��I�����\����s��F[P�# z���S6����p�B���������|����dN�x�v�݌eX��J̉�C3�ě79�GG��pm;��e"�����'��[�U8U6�o�;�t=#�}������ �Q�};g4T+N��c4O_��/�:ّD0����/�-��˯6��1<���d)#���[�ck�|����"FJ���
e�3�qͳf����+�VY�Ӆ%GH��g��`�
Q�9�X�ҹ��L&w�"�;�6�P�k�M���P"�{�߽ �0W�	zٝI�|Og?ݍ��h�1��F�>p�@O�5���V�;}:��0o&������){˞�"�.�{���bj�Xe��9/���1w?B�Ez@�NЉ
6^��:�w�!YR
�ߜTf�R�e�+sSVT|3���S�1ʺ�`�nzO_?`<��΃���m6��?�E�}�5�Oz}�{z�-uW���hImV�_]�샇ȝ��ll}O��E5�9�8�g(��G~~A����	�-�(�V)`p����g�JF��{�|�q��|�������� �YUP����yj�޹��4���^�=�u��{���ի�t�[*�^����� #��eru�p����ڞ��\�B?ZY&��e�〤ܧ�t��j�v���Z�$��_��Rq�WO��ߒ �*�����0��*E�K��!��WC{Q	��HO�-hlk]�5T�2���6���x��-��zl:KvkKü&}��c���D��s���C	��F�x��GU"C��P�M�t��8�Ҋ�N0oz���C:��7�?Aw��(qp �R*�8�
��=��{��:�r� ~���n��-�N�5��B	:N5Z�n�O�x���>����
��r�V/����б/�k_�G=N�`�"	��4,>��H��)���pg�K�ᲆ�����nx�@O~��>oί�_\#q�L>{|��kWA�����J>�䅘�V=���r�۵�+8���G��H����.�D;��cJ��i�&
S��>99���WA+��a�cn�ﾢe2��3�BX��&���Ҡ��L�ׯt8��w����� n��.��oh�=ǫӘ�F�$h0V-��+���������(�B��`qYgSh�}�<�����Bۭ%z"���bX=��������d�rL�%��);++fC��������PYM0�g���Ԛ+}����U=c7|IHH`��U-�wUȄGX�>=�8/qm���p��`�����&?U��[�oH?ϝ�h�Kx����uXP�ݛ��fu�f0���/%6��a&1 �C�ۆ��wmb����=��b�۳g�XAg_>h�dP�)W���e<�@�������܇G��S�s�����l���|��ys��f�%��mu [b�^�ŉ:~��i�?�ljk%bz�
j�,�֧�o	�:�֤�O���� 3a��Q��$\M�S$�D��[iXC��7><=����Y1ݭw�hi����Ʋ-ʷ*`�A��;�?xɶ�����8�3�7� K�B��+g�b�҅n6vK�!�<Py�Er��.Z�tg=�u��l�p��(cF479�ea�i��g�|B�<�����������I8<�B ����99�2��5��]�e��.�2��~���r^2BKӨ!��9��g�}|�8_����+]Q� ��9M��"�7���<Ck��t��FS3�j�ߔ������/$��30��x`����D
���<B�Z������V��Ʀ�{N�dC~�x���lgĄ���]P¯���u�E��Z�o�
�
�9��F{.�X��3V�1�׮d��v�eDr����1Ň�Pv�*����߽|T|u6E�_�gS�T�:��bz�(N������ɻ{S����7��-
�0f��y�l\-j��#wE�{�:�G+��;e��E �+Es>����_�䉗�ǿ(P�l	� �j�*�/=7`����o��z�R��S.:�r��Ux���_��`����%�����K	�)0W�w��W�g		GJ�}L��L�I��N� ��<��sf�� �[�R����qʅy�2e�劄F&��Om���eݮEQ���u�@����O���Q_�l�)
�g_����|MDv�to/�8�_�<�A��%8OM6���� i�k{y-��o���@��Z��n�?>;t�yFA4)���;㿛�5�~fa��ipgcj��:2�R?�B�(�Q ����������<=E��6=�B���)'�/ zSS_��e���oy�L6��A��3��Mn6���xD`Jny�'��Q�/g�d)��o���\��+����b�ws�y��H?`��AS.|n0#�NL<���bF��.��U��0��KY�Y�d����&�n���;2�!�r�����0[+4�*t�
+�W���\5�?� �c@+G	�e"�@z�XS}���1bڑ�7��<�-彺<t�9[S��$HyjQo�ɗ�.�x���K�.�>�@�0�����ou�0  �VlQplՙj=X-v.s12SW�Z��!9�!dj����o-@$�����A�=���ܞ���C����nM���p�m��Vg��/ˉ�_��Lp�����!R;Y#�ts�&� ,��m��JluT��AR�]�X�����3���/�	��ζ�P�3H��PeJ�uζ�ӧ�� k�,��	T�@zeL����%�B�Fg�[}"���)5���E���ȵd�� ��tY{�������MO�{(��)��H���C�f@�>���#�/�"�
�h?���"풠�5(,4;��b���Q���?�uI0�9LI�	����rGc��Z�$ ���%�E�S��bM��������=���>2���"45A�J�#J��Z6�\c+�Z�|��^��a6�7�9�Z��߀�zh�]��W�@�O�}����e`x��N�E�,���Hn`�:��.>�ɏm��UY�[7�.e��S&�U�a
l˘q�?b~�{���5�wiy�)��Z��'6���bbM;��^�?��m�{��C��o��K`{�t���$��q���'�o�y�E�Qgi�i���>�a�b7����5_EEf<>�Sлn�=��c�xmԠs�_��xn�Bg�����m��9��Tw����d�t�#����L���o3�(���SHTKds����s��o��n2�N(t4a���y�Rg���(�DAuOϦ��ԯ�l�J(]�@�zYII�T��O�f�"���^:���'H�� �����ҟ:O)W�%��0��J�+���/�"��ᩆ?y����U�(N�L���䤵��]�Ԁ��B�Ϋ�2�QU���N�n����
�CM1�nh�yʯ@LK*%:��w�J?+>8r8;]6��+̉���
],D�+~U�aץ��Tq'(}�2��sΗ��V�����E&�/%���HQ$0��3�2�0E����Z��߹�� Χ?>=���	G�� �^9����@A��T*���<�����[i��N}�ME��������ڋ�H�+����Yq9+�������Qg��7�rP/@B��WP� �K`"�D8��}��j2�'������cx�?G(s�%]��uF�m�߁��CPV�5(���F��4����y�w��Ґ���=�%i�^�Қ?��˨��aa�u��;#�����ө�6l��k_~b��o:���N��2��Kh�8;]!.��kW���<��&K����d��ol��Y������L��ZSb�'��F�2�h�����33)c�����|C��L
�o ]}V�q��M7l�����yk���o�yV�,M��Y�M�\X�4ppĭ;����]��� �m�!��*0����Q_G���a��E"��֕�}wm�����ė�f�X�oF����u�_g.��HLJ�P� 9n&��Omy��RJB�̳��Q����A���Sg{�C��#��A}Ǚ�>M��J(�e]��{�����;N��l�\c$�]��b��c�(��?դd��
��nݣ_?�1y{M)�F�^,��ʂ��K5~Ʀ�	�!���Q��$[+�E�e��x���*��n�	��T}iiJ-A����fg��o���/�N`>Gg�=���ӳ��g,Єfn�ZO~��o�}����? ���z�Зb�+N��Zx��`6ByIYR�?�p�� �h�P�4�/g�m�EJ%�.���<S03f�k�D�OG�q��򱎈���CS��/��xa�]���s"/�;<�<��6���fe�j��#1 �S�II�+�2�9A��z@�X��/yi��4j�p����NB�\��S�D��k��*� l[�߰���Ï`�e<ut�d��{g:<� ��UX;������'.[�I�K˿`���Vg'�ԖWQ�az�=�[\L���3��ou9�n�J��}`�_[vdH�7*���qw��k_�P����IM�{#��L���B�4ہ�˓NLe%^����W�-5������:vw�r�i�yA��.���{7�M�N���~�w�o�
p]������K��P_��|���6=�����s6?,����,ޚӰd����*-c���(rFZ���U���N�����ላP�)���0��!��rCX����1�(%G���g{D�����f�fF� ���F5rbH/Y}{��fcX��j(��x9�03�\��oL�?�g�ȭ��ѹ�ա�*���>����x�ԪE %�sfֲ��|c|�Է�&����HyӈN���>�ۖ㘺Øz��i�~�b"b[@p:3k�K+ ��JT�����wQ-2m�"���g�����9��g��F�G�����V<\�;�ʊ���H����Ր��'9-&\!���8�[�Ft�U0��D�}2�I�bc_�?�%w��7������%�W��!te�����Ý�`�}Tv��@�Kee"讞-�pn���F�q�Ag*��%���T��ѻ�%�z@�nq	%-����'r+�îO����8�X��Z44��7Xc`��ŉl��\��N�{ދ]�w2>1��wW �9����&&��Cx�!*����~�m.��=R `��=\�W*�j�}�c	��22����#&	���")�Fݵ7��� �0D+�������A(�)��"�������t���E���m�9�w,��$�:���#��M��i�y�4g�� �)�x���ra=� .\n���H�brr�]��:U���^.BMr�={��LD�'���֏��~��>���ںH�=�%^?C��U羺�J�J�4��X-o���&�-a�S^�qyG�r� o��U8(9ygz����t��A�<^�o+���~ �h� )�nV�����{z
WcҲI$@\>��&P�r�ZLlxF�w�30� Nr�E0@�Q��8/��3ߨ�_U�6�P}�ʊPO�'�c�$EEl[R�IG�Ԟ��\�G �	�M�0g~������tĒ��	3�4~�]��%T\�\[[BC�SQ�<� ]K��n�)/�
���5l�hT`m�?T�@ ��>�O����q���b'� ��Zv�#n�̌_F6E�H˪�~*x��߽a
�76|����� ���ٙ��+E��0��{==�w�J���B��6uc	o�;~��Y�蓰�ܜPK�nc=eO.8�n㮝��� �j�	�g��61q���S�Q�M޴q��Mx���*�W���. q���V���,��?����xy+�#Cԭ� R�3���ƹ�&'6c����a��Ҡz9َF��,-�����[��6������3u�Q~��Ri��:آL����a�3�D`�w���-���/�es�Os.F�YM�_��`�ژVJjjʮ�;�KX���U�X�y�EYVߨ��ӧ���`��~xϷ�"NGd��r��V;V��eώyf�,?�r�����jθgE�4��60h�ihX�˟Ů�<k��QSC%6P��ڴy����T{;�#�y���J�ӧm@�L�
�P%��h#GU���@C���^���(�+��x3��x F(�|g�D�&�;4�����Ol@�ژY, ���?����3{D�����+�!!F���Cz�m�L�8R�X3�ﱈ�_�'r�K�6N�q)<�efU༢�K��Oҙ P^�˜k����N��g� q�-��7of��Q^��{1���3����huqqs{r'R��T����5Wx��Bs�[8 J	��M������ǁ��Ύ�%���gϘ�n�L���VP~���W�+���U]�;�}=fqW��Q��Z��&���(-���-��"�#d�:[Բ�PR�J��l-?�VOF����t[�"��V�qY݀��D"'s��T۳A�>q}SS8� Gd�o���a�zS��c�D��NSS�Q-QSK��M54H����h(�e����햔:�QK��[�Y���.��Iʞ�rS��HK(-.ݨ���5� +��1eG%&����IK�{:��\]�+�?{uIw)X0��$�|Vt5/osK���+M��sdFq���sע� ��e9����d5��F霼��Rū#T��U����hb�ײӦ�aiU\\���s��C���q?ƿ8���1���-����)滛"=YY��2j��y��"��j�%ݜ.�3�'�4r��� ۝<DG++��gL��\]Ӑ�{��?�x�7�A� Ô��Êv�t�;;\H]��[�^_�������\�w7�ݽ;����I�y�($�8�ˠ��ǎ���Ϙ�q>�+���&�l�:u*W�ԁɅ)�XZ�Gӊ���hb�Y��zcs0�P���G";���8;�Vդ�[��Xpw���:���"]W�9����:a��yOC[Gf 0I�p��3�ᳳ."2ȧ�:Q@���x �'����H��+��&��1W���3L�'`�J�]*jmhx��7K\m���8��ZZ&����XYv�!�g��:�,]D�������C	�\��V��('�:zD��bz�l��j\VցD�DyR-6�jxT��zd�`��,�lm}��^dhh$�k?C�Smh����S���w����/7T�YE�r{*�? �a��:������i�.��z�N�LaF�P�Hg��?XGq����mxex:��%���33��x,�{u�<�R2]qeM�r��z����Q��E�`����"Q�V��4�/_�~��?���
����g�05��o=��ػ|p~ߺj�<�`L�����a_��z��Ƶ�f,��E<�%׿&����>�_$44(ܢ��1�T)��$�Dk4�X�.x$��Еb'|98��4�L'+��ϟ�%&�����$#������#� ϒC�ߟ�Խ(�0�s�r�h��W}�I�3�R{Ȯ��j���OK<b��	�'Z1�.�n�E3������!������|aAƊZ\xCOIT�p}UC?R������o��H����(T��#�m��}�T���i�W��1Pkt�"XMc��~���ʽE_{�*du��T؇��Fk7T׊1�ǖ�L�0}�ç�~��3��b�%{��!�,��yr�$�1����Su�u�U%��v����Y�o���}������*@�!<�jP��R�=���!�;!y���`F�o��նr�f�~=]��>�Y�c%�Q�bK��K�>���.��RD�t9�k�\��{�M4ΞF��<�H~�P鏉��h��k��Ϝ�z^���U���q:*Z\yچ�z�gzh{�C�[����޺�램��� ���i��y��**�����P�Oc�!��q)�{P}��>~��q�ܢ�U	�|��C����Đ&jB����w����.M�0�I|�9��b�[� [�gOk�/N8��p�v���`"�$D���҈�X�П[�Rƌ�ש #�?mja��]�j����@%]���߭�yP�g�3|�]+c�MA�A�ꡖ����iS����`��\�ę=�w�y��؏�*�T�u�Z�����U�ɑ���k��W�=����J��[���󈐀-���m�(�2�Z�x,�r���渹K
3����7�O�s�b�'-E�Yn(��|��_�ǵ�Ja��n��ǵH�i0��kt�JM�����
s����'��8�?[���k��v^��v������;������;������;�_������5	|�a�
���;��؏�[?�~l���E��ߏ���'�~l�����c��֏�[?�~l�����c��֏��/�.{,�����+�n���h�N\=�W�	׋1�1�
��xo&P�\���<TQ&Y�q"Ź/��ގMH��R�;iy��������˿~������N��O�Z�����1fj�]�4�-�+�k���L�a��I��]���n�B��������^�+���m���BߏS��������){]З�U�|�Y����7zz��꼨��Y��=�)�Yk��?}M�jk�a��S)B����s���������tA��*
}%���t�@õ�9�񋰽�,4):3B�*J`���B��e6�A��o6�o����k�.	��D���q}�������>���o��M����.n��+��8r�[�����.�yM���|�C�?<��}�qrq ��7��/�m
}�:n���̌��o�µ���T� C���IP�١\*4�ۥ��4�b���Ŧ�h�>��p�FA�����;ڧ�//]����tH.n����Q�O���E��[4:>�/�}ʇ�����@8��M�Pl��� �4�$������U�]�y�A߬p�ɑ����B�{JEK.�߾������LE	�7%lV7'����τKF�u�߰�y�;�d���z�ף㟣�V*q��/)��I��Z$��צ����C�B�����C���!�_@5���(W��(���v�Y���\��k��Y�i%�hx�r�?���e-V��S�8lv�\^t�W֣���|�.Q���#���@Ay�?v�e���VrBo�	�������YJ����Q~ڠz+Ep���;u%����;ڿI?��B�9q�M�+��4�O�(��ۂ�d�v71�g`�9H\Rcww��t����971��ndd$�C�o��7(+)q��⳱o�I��#��!VI��v%� ��1@����=�"**� d��e��"�ww=�+�]O��@�K�8��^�.P��f9tO�f�7�:W_,j�����C*����q����PY�}ee�%���;��u��e��OPS��0�L��6t�2�!�Ԋ�	�J�eqǑj�`��������M��	fbb�8)@P�p'��\�kI�G�D�8M]��4W�7�u-���� _[��g&*�nD�Z �С�Y��X��ᒀ��9o~$@K��S�FPj�7Pm��_�H��C��\X5�+�{�5�!ǵ1ƸlA`�����̲\TM��h�m�"�g ��`%��*����b��am)Z��ԑU��h;8�-类;��B��uG�T�J�`��1�a���v(��t|���V�'wwu%�(2QQ�	8x��M�]!��G��X�!��̃�ammmVV���Co~���  ��'Z���kӔp�ySllk?ӆ�?U�#᜸�?�`�M�---=�d���eg�/FO��srh�A'�?:�0=M�*��P�]�"� �ꈟ%09���T�R��M$w�|��&����C�$p��E�V�"�˰�K�vF�Z}O(V��ZN�е_ @z��J��<���~<�팘�~wR0d|G��ˍ�I���\�X�w��f`�SR�H�4�ae6iu� `���LNFX�p)B�q��8me�������ɷ}�`àOܭ�Oc����u�;ݎ^P�+{�1r�4����x��R�e=Dˮ��~@� R�;�ӑ�Km���ߎ�y�ǓQs�+�oBrr:2c���gԔ�$=�����-�.� *��/��P��Cm�8�����B���?c3����I��$��B���� T�6k
��Xv�@�P�^M�:m-.*�HPv��}�\Hs�A�ǀR��yH�� ;� ��"PR�R;:/�z�j�#��`o��	L�MR��?��p���S,����.F�r�p "�r�ɣc�b��b��N�-�'��GZ�w�h\T:�Z-�vy���G�V@E����)�wtv2�.1�j=�zn�)�/]����W�ĸ���v/{��2�̓71�����UU���j���l&EEyD�$�=B��� Q���#ge�+P2�1���=�	���Afi�8( �p��0P��%�Rڱt�g&���Ƶ�}TO���B郻��I�'��E8 ����mc8P�:7A��^��n~��ys�m�)Z�|R�yX��sH���K �� �')U:�<L��y��0��yj �C�2����b  K�{3)rEE��9!^8�r���k
gAX���J���f{ĕ_�컀�C}F����&��*�*�Y-�l�*�hY~mHNN>��Zh���#��azT��V`*ճS�h �E��������Ǭ�0Y��� y��׸pv@���U��tP��g:�JKcc#[F����815W]�CՏ��*F��h)����g�T�$��
���Gb�:v0�p`̗��!`�\>�.@����L���[���� <fa�<OL��֦X�q�[@�ٌ��1�Ud������Gd�����Ǘ�&
8n[����EnJ��{v�6���	ǌ2T���A��3ZUV��0>��z���<� .aąs��93:
A��:�D�޻�	�7T,��Mb�\\!vh�|��)��������J�j���R�`�TY�(Dl��\��@Ԋ"�첷V��P5
B ���,.,���1(����Md�fNr/���?��9sf��yfι7�l�w������..uW�Ӛ�Q/Q�����u
�4���yw����:��r&�OS�B�:K ZG�3	LC�c��(A%#�M�T�pG�a߻�fӰ�e{$�~[J$��эw34��'��\2�/�d�OԾޢ;]UXs�x7�j'��-�8a�!�w�}�V�ߕ���?e<;D^a�\汳��> ��j��3��O��`)��}�١�|9
j`��N��)���7��9@�f���`^yY����WhlM�&P��'C�jzw�H}9����w���9(�Jm�#>��&�߹��G�-	�-n�6֖���4=Id8��f�~��c� �u�x�<sΉ<mA�:K��[?ɉV������i�R,��5&���$�DSe�YIKe��1��`��u0�qǿÔ��2�!�q~u1����n�A�xa]�%�Yi���D(3uJ(���_��16�i^,�6��v!8�'�el��$?�)�QHXN"U���DW�#��Í(S0��[wz�����ˣE��d�4��Ӣ
=���O�}R��*�}q��I�o��(T���zZ��)�7���95������w�/ 
||�c�k�J�3���b3���p������R�c�w˥�͡��wi��T�cPo�|���`�zT��vH����x�wO.��n��2�ǒ������\qy���3�W!�m� �Rh����@�]~2eTT����0_*5���nB��[˲;��(p���~� ��c�_W �E*��E��2e�W���ڰ�
)��z�ѥ��̢i����
K&�<���v���nkg�%���\�%~i���B�&&��A�y�D��TŹ��սc�"CD��[�0
B�)O��o*�}U�ݺ������2)4*J��x,&L�qGam��/8�Z�6D�oPk�=��!���<y�$(f� f*z+D�����HR.g\����m� ��<�,0hEzMލ�ք�d��x�rf��4.Z�F~�K�+��H׼�81��]a�oE�v��G6����'L����e�T��>���N&�i�5����6*���h�y��w��#�^����.q6E�Zq�_ډY�݊�y����5�&[�����`-���_Q���k���E��]�Zρj��]��={��5$�S6�d9�o8�ϝ�s��z�m�?��pn%�ХH3뚛�k�<=,��>��R�c�����
=?��DD�{�מ���2p����)��@=^�y-��>ҁ��{��3(�����
[�M��y/�K��j�;P@�"������Ԯ�\�Ө^ZX5�t��"7���V�e�ye�l���?*T`�l�D�3���.R�� '�.T�3������_PK�C�{�Z5�{�H��gKK�W�P=�/�۸�8^������%zz��I�Ĩ��]�($_���8�Z�L�$��c���J����T�[ePA�W�-n����i���m�YMt��I_�@�h荨b��҇p~�ܨS��䘥�U6l����DS��!//��I��d�T�*�z�Qcwp�p'm,���-�I	�5�F�k;���v�Ռ�u�?�ZRS6t@��+��%}K̻��3�+"㙪�S���Kz� uv����A�l2�q�בV��<��dk��z9L�Z�
'�n�R���b�4�w� 1)��rp����gz=�?IzO�f�]o޼9XS]=C�`��=���C�1��B1M���׹��5\���'_w�b]o���I~5j�t׫��P��u�\ۼM��(USv�p��p��P:���{E�w�׉�r,�78<�y���i
����Q�\��&��+��`�IB�u�hx+���_�����eb9���'�QķG��wqr?cD��Hz>%:5�`�0���ҝ{�t}U�D~��7����	�gɦf*ԸK��Hw� ������_�>gK���^3a�u3v�,p�h'�x��J�H��aN���s���������lIp����)֥�pmF�E�����$4_Y�Xߒ���Ιk�Ԗ^?�e��`5[m�$��)ƊL�"�Ҁ�����89�e�y���X`kY
_>s�����'�Η�c��}6�}b� iU"�Rm¥�Ӈ7�Z��N��}�.ni�E.����[�,;�ߍ��]��<�c9�!�Y)��8�Y����$�h������H��K�4}iU�Y��@�tॏ��Y�9/�8l�x�m2�]���Q'0��V��?�1μ�>�A�;�dȰ,��H�i�ĸ�E��^l��
d����o=^��-�x��	n�O"�������M�F�6v籃�mR����(����!�W�T-f�3㵼��bK����))����E��%دcc	Z<uh5��"��\��s�=	<.��J�������C��į�Q�L���c�!���B��jL�w�<L������X�$��5+It*�����'��LU��� �P�4�P��T�"��������q��I��h�8ހ��c�C?Ț8P�
�$b�2���<�V��S:8z�'�u�H�l�_X�o_�4���?Y���{��s��7�gXֿ�b���{YE���߮NO[Z}��__��u��k�������W�t��/�}~�r=�.�L�c�qo+?�*è�Vm�ќ"���Qmc���_+@V���]O�
7��}���i��ɓ'�$�i�:EfO�BG�y5'�[���wg�tΘ8~�b�=.ەi�~X�g
�K�a<��d���p����P��WۮA��3���jhd[�#t��-;������{�"��[_<��\~��օ*eKa>�$�$"�G�)NH(8<?M�H>����4�./��H=���7���t�yc�#!hU�i�����[�N4?�w��؅n'zӷ��v�-;Ў�AP�w=7�KGy�)�����x����H.WhAƪ�(~����F	b�ɅB��O�#J^Ң�$���P��A�nQ�-�����"��ϧ۴���~���7�\S�Qk���ؒ��F[H�O�[�`w��fO��zG{ޥa�)�l|��Q�l5�竅D4�"
�{��ʤ��?p��W�,Y�`�<��1����\nQc�!ˍ�z57��-Mt�_O|w��rc�Н����"�kɳ8��������(T�⤶ƢQ?O�٤1[�}1��9b������L�|����������}~V���Jr��+[����-Q�J�vg%:i�#1cTQw1F����0��� gWȒ�---}iJB�_�mHN6fv>���gXT�co�=٩BgM�=�Bg������Z��l�AvM�y�ۤVG��p�� 2��w�L)'�b!q��J9�� /�]�h �y��
�z˥�ÞQg�ImO�Ԭ*QC��}:O�(A�+0��������M�J�f.�!L����O�0�ߝ�ȑ����*<����AuuujP�9X�^ÞQ�Gb=���h4����>cSJoa�S�2���B�z˪"�������lkW���6(�V��0�w�z�č|�ԙ�o�O':��)b6���8�F���-8L$��6ZV��SF��@Ss؇;d�>|�pgHȈ^�*��3��*���ǎ��Jf�������J���s">��(l�Bh��_�t���C��)$x�Q/�^7٤��m{�YfW����:v�<��==B؈���|�Z��|�L��,-3�B�p]DP.*�kw;���s �MzxyQ7�Т�Q(�F^�d�����k&�=�e���\[�����k���]ޕP��N��W�������G�[����j��A���+E��|���~X�@��8���L7�����ۥ0b�
��w����"Cm�w7T�I|~I��gݻ�Oij�Dyo�E��?�5�)�h>��kd2�������i�iɻ�H�xy�����s��
GmqQ�o@ na��� �L���_��u\xO��ΓJ,���y�u_����5f:��5nٝ�b��'!B�Pa4Al[CA [�s�l��GfĮR>j��(�0S�]͊E��ڥ >1-
�יe
�?5�w�fGp�ߨgv�It�%�,Up�����B#-�<t��s��?>o�w2g�H��82�/��v�^�E�Hff��$uá�D!O�R
٨�#���dN�	�yCh���a�}����F��J�1�F���y��Z�p��I�����W��[���۲��݇��B2�<#P�w���O���ų^!�v5F	��)�1���ʸĜ��ڀ��;�Mir�Z<1����������s��c����ξ��J���<(z�B��)M�1d�k��u��������I�tY��޼��?��#�>&�`^��"�����+dwhF��{�5(�-���P��{ o�II�ƶb� n�N�-�R7�����N�vVjʶ3P��L�(�Rw7B�@��G,�R��J��T�vR^ug���ѣ� ٜ��Go�Ȣ�޻w�Y�;��MwJ��4�b���No-O�wk�S�G�9����9�L�:/
s!���w�.�~Se�hNg~�)>�ȂL|�Ν;��z�6
�)��%��f5OA�S'7>��QFB�E���4.��aN�?q��?7��tM=� ����V/�	z��"~n~Zk
E0���@��R��F�w(Jk�����J�MP������)%S���i_�Oi#�`��	�2<��n��^���0ϙK_î/��zK�WG�2)
��C�ū#oƐ2G���3�����������\!�+A��S�%'��L).�ް�s[��nS:2<8:[�3�Lff �0�ܲ�����F�w83�u ܘ�%����Bn��u���Nl�
6Q*�I�n�r�װ��ԝ^�P��bD�R��?��s����� �`��@8|�[���(�LE֯3CGG��sFW��8��fܺ�Z1��}�@]� bX���G�{	s����2����K�9�(��F���{z��$x9�A�6�T��+n^�}���g4��9�k���Z	6�:���DR����{�i�&�,�Ǯ������|f�)�������J��k���v������hcJ/� ����:@ �qM6��" (Fg�X�{x=�ŏX�v9��
�b?S��� �L���H6�a2A@�,�&�b#��
)kZ���!r:�9���l^���j����H�#�Ϗ��n*�P�u�'��J&gj�������^	[C]��X ��|��<U&����D\s6���~M�dB���#�}ɑ%eն���4�6%Z��0џ)MR�?/��[E�*��O@/�k|�%��s)LW&)�Zka�ZY��j(�] �;qK�?G�l�k�!cѫ_���5���<�q5�)s���d�\��=��-�1��]MԼ��Q��\}�5x����P�&�υ�VO|�_N.��_'1�'?���X��iS~Dx�tt�b>� ����Eɕ-C��1JO}ww���aP�5Bé.]��z��l;;b��n`샱�7�֧��G=#�����A�Uٙ�oĝ��G�'&֢L|����Os��*�W��v[�:S[?���N݁����v54\�)T��ׄ)�������BC�@�����b�0����=SA��h/D��Ľ��Ə+�M�i���9����[&v��}x�#ۈ�ϙ/4�(hx!� GK�^�,��m��0�.��OtvvN�b�/�8%����]��,Gi������@_^�v"��555�j�N&%K�%_�O�$j����qI�R۞��Vc��d.��R�;(��i&%	�o���q��IwB43�Y-��MgFa	�g����N�9�	���$�a��
�F6sU�=�SZ�Ty�=���<�p�I~i�o{�n~"��P"JKk�t�`�EI�C����Z?��� _���?F����@F|��-��"�\'��%m����9��ߺu+��0��oi
�6B��_M�I $������3�~
A|rg�7mU�1~�����0\��$	�n�on��s���7 �����f�
ןFk�0��RB�pB-�٘āOıwRO	��P��%�%Vp���ɆҨ��ɅR��Br�^K�Fs���-�w׎�wS�;��-���4�73��)n�LOq�KS|�mo��#��"��%$aL�1>/J��k�����z䓡[G'����y���3�/����h���_-n�ĴM�9�52"�+�/���e�i�0G}[Pw���5iiD5v�(����p�h;G�4�o��rVH^Ւ�$X𲡸4!9��S�����i?�J>�`%�x�L\�:u���qS-Ε���m����>l�����Z�Qw2�����Y�a�"}��2Hm)��n_��If�C>m|-N @�! ��Yi�1o�[3)'���6�Ό���H�풉C��bn��(�S�l�6��ajL?�dS���s)9�m|�Mu�|��w�K;pQ,'I�=�ԩ!c܀���x���+[b�힦E k�@��Χ*�"�N�����3�� ls�dq~�o�U"�v<���z����e��L[u)��
�4骵�:�;sq�VNS���ýGz�e`��uF+;R��?inn����÷�l��M���JNA�i��Q����?��>5�y	?0Ց9,5���լc��fz���WEE�qS]����:�+��Bф��&YB��q��PU{�{�^o&k/���.�l	�͊��y���\�5#�$#h���a�?B���'��&�����Cjb���s
��7�=䌨�A"
 B�E[�Rq���l�N(�Ĕ�B�dh���S/<�Gaů��v�&�&p�t��"��N����fH/��	�R��g��<c��1��0DކA�̉��c�|�8����Y;8�ػw�I�w��Wf���5P!b�f�۽�L�V���B>o�O �lV��.�{kJUn�SL��>�C(8�@K�M����K枕h��-C���XE褛?�9k--[������b'��L YO����|K�р�C;%��$���$`�v5嚸z8u�A�Mm��{���=�nu�'�D�&%>`���J�����ԏ�;*��|Α�,6�$H��S4��{4iۤV[���	pxlY����|�xj�K���+��3ձ�W|�x����d+��r�gX��ˆ��a���/l�F���|�B���#�P�Bv}�p�����-O���[Ba�*;��0`��=���7�ŷRU�z�z��I��s
�W~:6yv��[0kͣr[��6�-9"o�0�z���:��G#���T[B�*��#�SZ>Y����s���K�b&�춃�Ozc�C?��N�h�pܫ��0rēA��a���6~ˌ�r�Ġ�;��GIc�4��Rq$��#B	z�K�J�^����
�d^�d��ifl��d�L=��tBXۨ����ͭҁ��Q	q� �J�u�]�B�kN����,rP��[�����I�O�h���M��`��/ ^>���֒0=H�bQ*p�]�-x�f�,�+�®F����dj�D��3�v������π�+��Y�=�{�����D�3=�5��B&�\Q�	�>��$ޮd�O�J2�b��iK�o�,�N��e�}�W�)7W���g����)��׵���kB�4f�x���.���$'_��Ѳ�^�{um�y}�:�J���F�P=hM/*�CS�S�|}��1,��+��m�"Ɂl�×�@�mL1@[&xI�I:O��n{zE�Y}C]�9��j�������li�7/؈�?a��[��=X��G�)t�*����#$J>�"��/هz�C�����.y���7�=]�3�ض�\i�W߫B:Ŷ� 5��8�oyb�l�7T6YY�[#��_Lɲ�wa���1#��~�z4��#k�/�B�%�Λ������P@�`:��sێ���9�U�h-��
�f*��s���PX�Z?��P����ɌMh��$�K.�����'��bz�zrO0/ �]�vͮ�g8H���b-�#h�˩�P<�dسK7w/���J���U��!���+kb?���\�$"h�h
)�.{��9_�^8��K����9w�x}�����O���̓�-�P�7��}Y6��V�6��7�~��w�p��`�Q�<9��IĤ��$�PW~��ݯ
�g�G�>���H�ܑ�hg
~�+�k��2�&���[�6��_a�ap��S[':n|>�M�-oFۙ��"Uf	j�WB�8�cJ�L����kZ3��1��A2�2�s�W� �� 6�z�fiE�͉��e��,�#_a����Ȏh4�N����ѣ��e�T���%�=�0�ҕzK�4,V��N���)�b+��D�W>^�ũ	ƪ����xH��	
n,���xw&Q��l�B�F#��^���-P�O��oM��.�+�ܕi�.R�I؃�t�;�%�$Bu�����YR�^�2�О���@wz���!��<{�<v��t������.n
��G
��^r��cK�ÅE0-�	����Q��Q���i_vm�\��0z<�����9��&`�{Xe/SSSup�u��XA�%�ʕ.{4��e�)���eo�ī2���{�ؾ�e=D���)�	M�zܡl�[U�.ǀ	^=�T�|� �eS
�s�@��	�1�N��ìq�:��-Abc�z#�jv�������y~E;!�_Dl�S'a__��WS]=U���\������hkkc�Ǒ����d�Fë�]�H�+��>|X�Qei�0�����M�Q #S,�m�YV�n�,��Fq�[�O�5ڃ-�k��zȩ���y���^��:Z[@��wߔ/_�ͫ��O�շQ�c�ՓwI�yC�ȼB>#�w�<�传�w��)j�ͻ-����\���u��B���������P��W���R��F���?��7Ae�h�����%}p�ZM�Pi�Sւa���k8, ��z��*K���Hl�-1F����Ta������*���-`�y�M�x���vÅ����n�\y�'�ƿ�fa?^�~����]=��d*���rb�k&8�W2܁>gsK�L�y(&ѩ0��6����x�O^���d�t@�s<���1�5BuY��E�q)�k��=d�z�F(0�:
�I���@'?逦��9qѣW����y��m�+�H��)�,f�6	fv�S�Q��ᐢ�G���;�r���[4(^����I��9N�3|���f�1���+�1^l��[�W_U����vZ��-.NW�{%Wzi-k��+����J�&W�������w�)}{c���7_ٝ]�W��{��O|��-��EM����}�hZ[�Z�� ��s����t�\.׮�[2ͤ��s�{kϑ�iji��`�\B��#��o^Q�W�/W��)��y�!�(��H�F�Pb��MK7g/�	�/�a�pϓ'Oҁ�����ȣ!r��h����;{P}���ȘD��s����p���	}�;SzX�M6)n���É�NY$0�Rm�b�w�K��U.�.�����e���?c�|P͔�Xwi``������e�
bŃ��-�Z����@)�Ng�2���:����x"f���h�$�Ň(�k���ů�n�['�����Ǐ��kɄ�+T3�&A�>'�"}�`�̾�q�
3��2J9�s�]���cW4O�O�n��_��;��e"�gZw%i���Dۈ����I�j��"�Gݻܐ�esYD�K��| R�%�vQ�����Oâ���l��}7��?��G��O�v"� ���2�HF���ħnj��r�Dۇ�Qq�8�b����O3���;���԰%���,����LOK3��e���a����m�ήtw�qLF��2����C^O2)9H��y:>�p�L��dq;Հ��,�K��ˏ
�m�%!�+CE���)�\l���7�K�d���%IhMJ��2��$nn��+/�t�nS�D�	��}��>*�VBIfWc�m��B�y�l�}��~�ŒU��V�/V3�S�-���� F,'��+z�KK&F�B�m�<R�dxܺ'��(��"lD�o�*�qb|���
���hk��0�]��Y��`K��ml�#��Oe�L ��Ni� 2��/���ܼ��ſS�L���Ȇ��
���6�5�N�!kS������r[�*Q'�t���Z{?�5��R�{Xx�I~n>��gI�U���s�2t+�q�J�}n��Lt%F�P迣�1t����-+%����<�y��$x��0i���GK��a�l�_���WX�S�Mg[�`���i�]nJ�Y+ Ch%gѻ�D���C�&n��m��^.7������G�Oa`�[H�χ��vNR7��So�g�����*�l�ӣu��q/�̸� #�Y��{� �ߡ�7��ٴ��,�Ƒ�
gt�o@w�
&,Iu1�w���l��nZ�2_��A�"�!�|�:|>�FZ�IO��Z�~�?N��`�D�5֎�9�k1[��(*�>��/u��z�@+����Q���n}�h���Vd/ɢ�un�S�+����]E�q��k��a�k����bE-c�>L�:���t5;�:���^�w��<O�+�% ��Vd�c��7#}Q���R�Q5���o�BI�s�͔�!�v��ck"�1�-�v�q̬lɟ)���U��)�8�t���Üv�.��	~���s�4�[(����Ȳ;��t`DV֤�NMN1`�Og� gvF)=5UmW��)�՘��v����}w�Kj�
�x�tt<�r���Vt��	�Tb�&)su�<���D{���K�F0�"/)9�|^�	��2�f"��b��K�y�F��~|�~Qs��3tJw�z2�1E"Ga�V�/:J��PJd!�'��#E,��hG��!�~�Q�;������ %=8��\�%����*��VI�WVV��e�b*&	���շzJ�qK���Gijj.?�@�M��UM�mj�T\�d�[6�@���u3��"B�ڤ��)))I�J���%�Pe����=��:�g:�%x��w�����
�������ȓ(#���p���%
/5V����B�ק�R<y�^:
x�^�^���I�m�=[F]���֚{�3�	h��Sj
�.�*����)�0�XZB�;:��W��;���FԞj��6Z�6�|�}A�É��e��>�a�ǁ�����c�y�6�r{�n�ڥ-�)MR�E�C7��bF렶�𒪓�No�7^P��_�9#�!�~������Os}Z�k��v�� ����_�񸮮�!đ(/�o��Rw���WD�\G �����(�{�����[f�~/��^i�Mu-MMW���朲޲j��c�)�i� ���N>/����m��U��f�1�'�$j�K�4q�*c��`��-{�9I�I��ʀ R��O�}*�����KU�լ�lY���D�~OX�㟢�x�,--���s���~�U�kA��L�7C
��c{m�i~�w��Cn!)r	�8��gϞe��>����b9��r�,�Zc�Q�̶�/�Z�������﬑XV	3Y;��ބ\`�)�iRRC,x��S�w�1If�P Ly�3| ����@n/������xe���)�>���ݭ�]Ky��ƺ�ӧ�Y vz�W���
	9A�P#�A�Ѓ9@��{h���-tڱ��}�,����&n�ٚ�zrp1�����z_Z�U%R����I�ۏI<����]���LN�eItU�1;����ӧ7/@���%�I�}Nh&����hIͰ�*���?�5O\`h;�	�6����>��C���_p����H����*=���Oڢ�=\h5�x��	�?�*Lw�J���A����"�ҳ��һ��W�T�tu��s��/�<�����7�dK��d^����x��{�t�$�^J)Z��"2eK���Iyâv���T��G�����w�"��
ɥp�r DiG%[x���	��O�~*�％��qhѐ�~�wL#I&6�I��D��H�֯�Z��^����+>��wEid��̖���u��o�V_I�Ç�u-��'��.x�J\�?$3m$'�c#��W ����=�'3����99����t���PM�s�|�l$��͆-il�0�r/̖�ʲ*��yVs7"��^��4����YjH���8 ��!KEa�P�g>/��oP/�QeQ��+�}*���k#兑�,�����[�v3�m��r�����z��t���ׯ-�΢_�=�)�*9�>ګA�y��U����2���R�S�̄R�6�Bq��/q�94�ï�,�����2�ZEC�1,�ܧ�*�RgSJ�EaN!�W9�=i_�H@��tG�ֻ%Le����J�`o?��h9QJ�`N	�i^ҝ�J�s'�x��63���>v�סd����GF���'KD!EN1��:A�9e�e,-X�vr'��`�yqwh���N��tzN��v��1G�+Q'6H�Z��\ûh�ik}]�������*�Ϋ�o�B�v�B��sꀗ%L��I�\h�*���ak��Xc� J-̮�dM@�*�}��N�^e|�d�Z-,,d�_�Η,�0��:Ρ�	u����T�U�,�ws\���Ȩ���5>�D�Ә&D%ǒ(Y���dVٵs���wĹ���)
-"ϓ��Y	&�jw��@�>��Py��%$��]�~ɕ-A��݌�ɆHo�����.ج�!�zD�����Ѕ����{}p�y��ڝX��N7�����5����<�/٩G�M��dD�K�������/�|a=x�z>,A��l����g2י���ٳb��-��lTH���SKK�#�J�frV��\[H�D��MU�!i��nj��>[>�LM��Ԇ*�Ϲ*[��|�ߊ����{�����0_J��/����T[ufƆy�� \���3L`G�a�o��)Yr�oPt�`��=�r,0��ݳX��%g0.8>�}(�����n���z9/99M(L2)!��rU}yP��+�.i3f%'xI�T@�ܷ�0xP:K9L��9���ٵ�2�S��䔴rGw���*�cդiH.�>���~�.* ��H�FtI�����p�KLyN2p>'t�C�tl��j����z���NU��ʽk���G:�y�ƭd�B��K�C�� +}e�Q~FqbL\�]J��Y=�)���uq��9���4���eW=QDV2��jM۬-���cc���I�3�5	C���Y��S����ROi�Ye���ߌD�1���H��}"u�8���<�L�*)'3��(������ u��������ڎ�`�r��kkk��� �J�~�Q�qdA�x-�ɰ��:��n!MT܁c���������wB}�k�)Bs"�͂���^����ID�$Ok\�l^R�&;@���Ν5`�	�RR/����ͫ�F@Ѥ)��Iy�~e��*��%���3lQ�ѴvW�''�g57c{��)�7���83q-�l0�Q��F3�ڇ����Oi��p婴����swϴ���d�>/��Z��ݘ��ԡ#�1/�r`W��:2�:��ws�-�����Ɇ��X����[�D�Z��*�0����y�Gp�+�4��$=�)���~�����$B�3�eH�B������0Ԝ�M��B��k2�$�g�^fW!�Q�	>S��m���W�W� ��$>������>hb(O0�T%��%��=�3�����Ɛ�hC]Yh`�������4�)��|���m��Ii����E���yk��U���Y��H���=<ğ������yb��B�B�y�-�B�ZF��O~V��Q������*!'�w�} Q��	ޑ�1w��jFX3ԙ�İ�eG>��χ����C>ݝ	�E7�zDT�u��3[�H�b>R�
��1w�¶?Z�n���#��C��v���N^#���X�pA����:{�厴��6.IB��$:����<�L�Z6�'��i\B�K�JB]�,�jL�8|N56�@A���Ax����=��s݇��cS���k;��6YY��Z ��������0-Z�og��Cq7��k�Uq(�W�nT2f���۽���̮,����6�m؝�F�r�=�T���aNJlݟ�`H5��*�s�y��h(�F�Q���PP@����C?��MOi�۾����u���f�c[Yf.�5�A������G��<�~��߹��(��Ogs�sds555��Si4����M��i"��6)M��(����? a��0�lo����vt����|`6-�R����*TT��,h��C�v@��1�Iku&w�|�ip((�&��)t0��$�k�%���la�k�Î��K�2�W{�)&R=|e.xρc�e#�===��(k��u��o^(������tP����g||�?�kqT�}ܒ��m��Vp�����TQ�T_''�+g5�[�3Y�{����E�_�*cRr�&����%�r�ȧւ�I�p:���\��x?��Ǘ���u��yG��)~�牀y��<z,7��]W�����5"}|W���ں�-��*��[8�����5�3¿�;A1j<�ѱ��E����i>��k�tP�!�ʀ�.���Ӷ����������	M�
1ëX_��ЗDlkC�V�rZkQ����D���'���ebL_����7_oY5��܆���4��4<���� �Y��s:���]�K������k��o�U�Yv4B��ni��յ�1ޯs9�)%31<6b��&�.A�}�%i4����W�2M�NF��P��台�X�l�jV%<`�Ѡ?���<��s�Zn���������~�� ]�{1��hZjj�Ld:�٢��-!�����������|��BE2����3Sa:�!�z�z8�³5�E,��+l:���#H=:�IkzVe�福��x
���$Q�r|55�;��
�Hm�x�q���K��k̝�?GL�f��>w)?��95c٢E�9-�^6/BM}���e��w�Io��~~>��\M���KC\�٧n��8�=����e#������"��y�17 ?�_�~���5{y0p�'�4��q4$P�8�T�ꄃ�z�S�>���_C�p�t���t�UL�M<�3�Y�����.7�sFX_��liiI:1vj�P�`i�wb�1��<��kZ��C�w�eU��R|�Ӈnc�<A7�%>y�)��n�XOybH�����;+�j ��!��VA�jYN�����'>�\�s����Pt�c�6Ӣ�Xȷ��w{�\(�/�c\;(c������ҒٕZ,��;�[�0��G�%��D����OvgگǗw��*�~�)��p�_��[�C��*@&4��ݧ�A'�sbbb����k�ل�ߣ�`��i�.BhD|��h���#,�Ǝp�ִxO277_>�e��EY�#kO�������M��u�bSB&6�'#���R���TIg,[�Ty��ah|g?�2��HGG|�_�	���R|������ii�Ȳu8��昁ǂ��d5�8a/��!��8vj\�f�(l\mB/\��D�pb h��}�FwH�0��i���I������,�i�6!'�=_6dj^9��>D��YNn��<IO�P�@�d�ڬv쀎P3f��w�(p��jw��V���� �GֶۓN�8��Z��
�N�;��sxJ��'k%���C!k
�iI<�ÿ8��
8�n�R��ͫ��w���&%����%�˿7A�Pv�14�����/�{����IY�m[��U:�z�����7���w1Wk�¬�*,v�W�ε́g�.T8F}}�3%�~�u�p�x�������C���Z�̼��;�����㠾�Gy�95����/;��[��������~�e�n]@��4�j�������/�yٵ����y��w�ZeK�6��UP�?t�/޾;�MD"m�0'Z�~�e����T}����.�Y�Ź`kF)Xm��m��i]��+&q@��9�e'h+������u���RO�0��u��.W,`�^4z7fgg�U��U�h�=���7>�	�`%>�d�ȝ��3Fq3�M��Í��N��6�1�*������hS��-�;=.B��;�ᒖ���{��~�Ȱ���3��Uf�q�ƫ�� ���`�4%	���]����3)QB9U3�����E��U�����/��̄2�	K�k^�����J�^v��4v-`�h�U*��^i���������ސ��O�mS�7i���Zң2�!�ʀ�>�h6��XD����6��a=�m[�M��+��o�{��jq6�d�͓~���A�f�k���\Xi�3p�!����ͻ#lZ;w�nu_?y��4G��t��X���F��3�.=۟}���V�����������*��*S_%�N#�}�����b�椇�!b�:>X$�]n��BՋ]���O��j��Q�K��c�M�zt0�T�l$Ҧ5��u�[���6f���G���ܒg�yq~SOK����.J�����z�P�F�rS��G_Jtj���`�d�����=@�0��wcn�8����`�����������?�e������%��x�J�q}�����\�2���k�x5�����=zT	�vqfu:*e0���U�Ɛ�������$�V�msO���	'q��1�L�Y��q��98�σ�jD����.�\�>m]�N(�+JF� �ռ�|�&5�w�ɘ��$O $Xp�tA��]�9�y	�(}7��t���eqkC٬B�e��i;��;�f����O���'pDy���=�ڷz{{�U�8�1+�· |d�`Ct
;�OdV7��"D���\z��Q�"ufgq��8�;�sW����{%��;AxYz�n�D�hl'��lݠ|~vC�U�7*�N�]��a�>�	***�?;����^���8�C�|���q���� zm���D�pH�\ߣ���.u�Cv諎��`ȓ�ޏ!3�޸�C׼��@��^oe��W1��(�,�ruu���ه./{u�$rF�H�(��A�p�?2�ќa�xJ��$"D�X\��S�|E䩈�w��[���骯rA����}��T����	c���.g5'\���ާ��
MTO7���G��S{�1����<|�O�l����
Kޫ�k�%QWQ��?������z��6_���6Z��f����^Wm�.��ϸ$�0�W�W0�L��,����2��U��M7 ���0���ᶝ���(������#�~c���w#��N-��t�B)��>zl��ߦdV+|�	 �i,�f<8���16���in�4@�ر�o�x?�95���-�	�f��9F�o������r�����94�O����<Y��x���O���-2�s�DdeR�n~j3����3�gc������4�䬉z��I�Y�ٍ���+ �TU&�s�H�=�L�\k��C-�u	(ƻ�g׬vB֮�>����O^UrH����ga;����G!��5K�S���Ts\����ɘ�\:j|>{U	�����o��i���'�]7p�X����x1��}��DoFd6>�"�:��Ym��c��gli=�dA7zbSp�~b�@�?�[����#��A#l��;�c�)
����xP��7����������z�֟#��h��	�:8�zn�����D� зy1�{�ٯp#g,��G�ؙ5����>���,��������ɘq����5�\n���s?K�V����$�1�7�YѰ�	x��`Z���s`\~�J��
~��e��_<ϊ�P�pD��L��^���7:�}6�Ψ�ǐ2\koCX�G��3��q�)��<H�S�F�ӈ"�0�K���K�
g�F~�k��~AO��?�Ҍ��3	q�Ol�I�9&�E��zzf,�1ow������Tvz���|�Ljc_�ZQ�Uy��1B�y ��Ŗ����/�G�u�� -�<�ƿ���
�h�$hث�G�Z�p$��{F���f߂�۪���-��?�G �+[R4�ŀ�u�vw���
Cz��J����Z�|M�����6sA�����1��c8�~�ͬv�$��,�d�1�:�N��Ł�݉՟� ��Km�n�<���  �MA�jL(��:�kٯ3�`Q�}�$豵U�t0�rf!��g]��hn�]���e�^^�k0Fi��}�km|jf�23ҟ�R���FC=��3�V-C�+R"2@�� b�Y�����j��]}8n=����ZSX�k��[�� <�-^�������C�;�7��hGe������2t4vJ�{�l͂�-E�:%���ڬ�˙��� �܋�˔�}J��.����?u�do�������K�@9g�����c[
wuqY��Đ�y~}�������p��Q�;��g�%��w2+>�����ID����&m�?��\q������\2�?�e?����ask�����7}�q|���wà��N��C�l��683����C�cf��R;�p��~�
%ج��+*b*�Иd&[���{�p������|ļ��`�TYc�}����/[veuM���`?��K��s�7�﷏�.8��ӳ!"ݣ�C�ZV�Ǔ�R5P�߯�C��׎��rvn���}9�.��xJ�ec��
�֔�ŀ�]�n��P
��ql�Ū�� /w#^%6)h߅���fm�;+�,�� 1c죌ǻ�Cٯ�A&����g?����@��6_��v�7��vt.���k�y-���L$���%	Z�;�4�/=�(=���^�j:S�I\phX�}%���%��5��r�~��� PK   SH�X$�8�l  �  /   images/aa130aff-16e6-4627-9689-819d55b5861f.png�YUL
��Xq-EY܊����K���a�RtY�_����;��kq}����M2s�9�L2�3�/Z��X�XHHH��Jr�h��[0��Ÿxl���d������?�m����p���d��e�j�����e������ي���&�D�	�F_YN����3�z����k����Ԏ����(�Gǳ��R��7���c�JMNf������a�\w��{�I���kD�b�K@�)u+h��,?I9=̚;�����[�(6-�r�d��CGG�%��+��1A������G �����B���	�A�eF,M��Lo���k�=�8%_<�3��5���K4�AlaA��~��V����6�~nU���٤�:Ƌ]��d*
����W��CMy(%.KL�)�U~3"`��&���Y�t t�I� �Be���qkP��r�<f|0$L(��-+_�a�� m���$�J&�a���%���}$?�}}����4��ۏ��˜
|<gX��m�/���&�f27��+F�lȏf�{L�4d
�"��)"eN��_���`��N� �W��ܥ��d
ڵ��Ϳ:��-�^���X*�^�☈"G��oւ��^���i2���n	�ii��}I� ��M�L_�n
k|��g�^�D���Fg�Y�U��'�Ԥ��������$k_{���A��G�1�F\���uGLvaf��<V��W��f^���2=Wt���\C<�m&�	@�Z�O���g4��͆R����թ�#�7�Ȇ�A&��f�vf5
�"����0��hż_�z�@o*���I�3Mu�l#�c
���H�Z�I�C3n���6���ﴪ�	�,�@_�7���E_��~��ܫ�[&�N4�X��������'I��^��D��;�d C�uI'��;�����L��ږ��!�@7�<�^�����	�ʉ��!Zv�pt6�L(�QbG���Y��XHZ�e�<Z�L�$��K�V�jN]��{��i[E3<ӿ����R¼�`�ӡs@^��pv�Z�#�A��4d!~�D��޳%�{����i)�*7�CՐ��\,��{�_{A���>�Mu]hm�w�bD!�$_`�12Ő�Y�D	�,��&���W;��uo��oX���N��������c����`j������{���c�sH8�0'ޠ<C�ȲL�Q�ۗy�ߡ`��#��Q� ��y��IX��L�J�{�X3�̓0�1�|'��f�9�CC�U{�'T�K�c0�W�&O�BMJ�7&�꠰l�j��������X.7��k���leY#zu9`�4;��w�}U�@�l�`V�[�Zl|D`�eJm�c嶚��lnQ|l��;�l-��|�8�Z�-b�P˪W3��OIƭq�:��KS��d�iؤ�)��)hDסQ����UU��e�K��iKR��@�^9���� ���7G��*�p6�����Ir����1�q3��	
�Fl�I�=m�h	� }9!��m�W�:�1�jC�����w�(��b�������l7��2�~xJ�֛}���F\��w.5��ߔ�h)UV|il��;��cL�{K��ty��{ �``���C��p�w�kz�����I��g�'y�h=;�@�D�{:j^.�m⅊��|Ǚ9����;R�ȍ�� 3����xw\���CTl�y�,u�v�e����Y�(Tc4@X�l?��%:��v�M�(��� 8�TZ6�[��_��Rz�#�E)��i�{�5��.�X�uj}\m�w��~&�e/���H�8���Q�/���H�R��5���_�5�q��i�V��;���~�++�9Q����9=�CK�;G�T�N��㥲b�=;�p��>�3���W��.1���E�����|��Kv4/�t��XTJ��6�u{��%Ǻҟ.���G@���:� ��y%��
��E�N7(�� 2�-���]�H���Z�  O3�*韭�<m\�����t�pz�#�����Ց��Um���C�nĮ�$�e����uesM�����?����pc"a�4u�hi� L���(|�ϯI�L� f'�E"��*٩��ծ� 9�-]�]�������S�;iSKn`Uȏ�=����R��8�b�96K�A�E8�կD�h�⢛ns�/4��b�#5���6�R^&h`�j�y�9w�T��ێ�Gy�x˞�iz
z箹�c�*�_�9��Rg��U]���,.V�m
g�H ��rK[}����цQ�I��X�H�����rZ�y~ 
�6M��
򗢧���A7��!ܡ1�@��I�ĩ`!�j}���%h�	Hm=M��ğ2�2���I	��F��[�!�Myv�LE)v��� 3���>�xj�+�Ҹ��_��a^�h�$�ՖL����q�Rf�.��� ~D��O(h7G#�<qF�[)�������k�mFG7fL�o��k�1ջK����r�W��o���2Q	-��k�z�Phiѕ��"0����u��{���blRxk\�SK�.wFM=gx�)���;��(DCR���=���}���ST�P؜f���M��9M��X��Jlָ�.�1Bf�b�^�����g���H��(�_��_���	�F�(�P��}�y�&(�$՜D�Կ!u�y����e��a��,2�R;���ٯ��=����"3[	���6�rm�E?\L#vO0Q�3g��ˁ��m93X��GS�=]��F7/�=6��z�|�y��0�7�#�����7�}m���4t��`���H�袟���P�N�ɖ��{[���4xʨaO�K3\�qd`��R��sL$����;QE�I��G)o�LQ�uz+v׺,��L��X����%�\��p34p��Ѩ5 �j��Z��g�<6�^ܘ��岓d$^I�@//�!R}�V2qPN��H��b5~�q�@ ��>Jɒ��3��?9��yb�Yř��s���1]%���Pf���&O��O�X�����S���cܹlb��Ya��@E>��7X>�J,#�В��s�*.i�JeyL�P��N���	�@׾q��/"�M�))��u�:�����T؃ZV&���b��(��h5�]�+��9��0�Y`/��|�~�<�����d+�_?{����@�U��bꎘ�״$�P�`oP��R`]���;1�9<P���Ιd��`��rCF"���\ջ�(d>�M%DiJ+(63�Cb|"&��x�xL2%ѼZ����CV(�(�aW`��m��R�E�o�j�SX�r$�h�cz@�S��.������/���kW��z��[���z�K[�tK�f(��z�ôڛ�I�����r��,�*$��;$�|�q���zw���ǜMh =J�"2�Ƥ7���"Q6�˪]p̻�Aզ�s��:�C����w�5�hxa8B�L��n{�?���(�͸nu�$��Lt�z-=
>�EO��M� =�=�pΆ�0٠��Q��e�Q����_����h9>�Q�?O$W�d��/?-��uh�4���)(v�Uh��CJ���/Y+���<�!�Uw�~]PP�����Qǟ:�Ǟu��o0��|j�sv�%�U�d16͉-���Ze��Z�PR�_Y���7�������}���؆X����Q�������)6�	��N*.)>�.�G{��3�L^�u��p)��ÔA�Q��yM����Vp,}(Ll�xh�����---l�PT�ruru�ޥ2c:��n.1�N�\�4�M��3�ť�N,��f�e�����5i�@�Aɭ�-YQ�S���fƎz�
�*w�ÌO�ƪ�����'�J�/���#�%��.���U/��G�+;�ET|VP8�FBM����k�WY"���>ފ�]Rl2�T'�w���QK~���O���҃��b�15fBv���tA��g�q�<QӳRolև̅����A�D�.`7����B���*��R��$�ka]|o[d��J�=Q7�FbnO��I7#b�F���3�|�T�#1��D:��/MV�u��Be������u8T��'�&*�c��/C��̊�|b���,5|%���l�W�d�_���V�{������)���y��4C�dZ s���NX9�[T�W�⍪��ѵ� �"*SPÅ+W!��q#���[Z?��Vl���{�w���	�h�i6�XJ�/��I�\#�)짎��~��x����@�'^�u�! "F}���P�����@f�kM���������`mO��3���((��MƠ5g������본��N��_�b�mjВ��W�O�٩�7W�}I�.N���وa�lF���ʔG���N�$so��]�S�ee���=~뤶��@��N�z�5��:�s���ĕ����R���5֣o���laӗ0���>��^q�������3��2��R�7�$�;;M,ˈ����B�������`��W�p\4�\�qH��� `����1�T)!ؒ�Ak�J��b]��%{���DW$����~ս��F`(��ÑuCg��F�(�+g}}��'��- A��x���6����n���#<�]��a�������{�c��J�,�5�p��qp#��R�ZX�S�/.t�Zr�]A��a�N�(6���_km�mR�c$�<Qq��)~�+���f�Z*pk��Z�f�͞Ff�/eꝻ!Z�@�`ḋ,����?)�*��(�<E"�3/���"���"��o�{�RX�N��/�a��ZU���xm��iX21�:1}�,aS缈M�rwg�xM�u��k�Ѯ��e�k��V���S�Y2�֯�Tw������o���];��nf�/��ŧ�A��\��W�o�@��sފ�H�#��3��m��{"�E�Ӛ�G_�U�]��K�i�,�E���6��tl��$N�J�%9��{�P#6��䓏�#��.�^YSx��WBI���7m��O99.UϹ~!�t������	�[z~� SX]�"{��#���7��4w�M��z���$�o�,lM��u�D�Q���=429~� �����AŚ��Zo�Fc|��a>Bz��
?�.j}�"�F�4�'OdZ-�QB����j�IF���{$��dֵ~�l�EV&y�˩ XXy��DJ��c��_(}��s�T��Ҕ��[��D����Mfod��%������Y��cZ\���$�1�\�Tgp�ڊ��-��I��*p8�C��k��Sm6\�������<� qN�&,&L��0���=��M*�+Nol�X�V�ډ���b΂��z�o�����ӭ�������YĶ��U$��H��)�5�:eW���Z���<��c&j�0�b�m�վ�s���X�O�0!R+"����U%���a��b)�[����z5g��x�$����Ke�����d�@HN����c�܂ח��):__8�$���8�+�Y����JG�짽�4�E�^y��5p\���h��VU٥���h�븏����|��^����ЉO�I5'�V�t=`�},R*G���8Z�]��Bg�X8�F!�E�����t���2;ę����+ݘ�V��L�Cc}����)[�-�� .KfwG���<8^h@`!;��6ͮΒ��z�Z�%݆W�Z>;�[��#���0�%�o~���<;z5D�)a-��X߼}��U����[��̸��W>[��
���D&yY��~�}���cx�3��Ey�1�VC����wv�Ӝ�)1���Ⱦ��L=���V}8�LRo��N� <���5���w��x�4����O�߆��Hc���]H�Z	Qi�{�������ɳG�լٲJ�����̸�V4�$E�2�z�5�|�R�$5R�a�qL�qe��"V������X��	�y_6�IG�41��n����@l"�oz�i�v�ɤ��KlP�*$La��B��g4��i��/��<�:�\]/����d�!`7��k��J�AVf�����Pmܠm�g\|����"݇�P�B�?� �jdԇ�-�#u=
n��m9/.��\����\�]��g5<�����y4�#F��C!;I�@&0S#��T}���wd�@C��{�K�H1��7��,���M/�K>���-N<�6��"�wqN�5���s)��G�q*%���9L�Q��0�wk��w���x>0.A$���-�?�˙6/�PDH���>��2�P����Eiap�13.�U�Yz�C�)|�s�VkV����#(V�ʹK7�������ߗ3S��n��?�p���gҏ8��Bقo�'j���BbZ�%��M;#w�"�⮣c5~���/��IseIu�/�}�m14ƷS��b�#�<��k"Vj�͇�[���V�o묆I��?DoA	�Sv��&��������d�~����6��v��h��=�X�?mΜ��k{�����6�c���W�L}c�w�.�S�~�Y�s�_ٴF�u��;��8���g�����QT�0�ap2�;Z�1''����>���˵X�D�%!�$�ʽc��V�/&^+lB��IJ�(��y;����+<���V�ܮ����z���Evu:��2����=���!�K�[�xWK
�il�����qn��>I���-��UI�rub�j�=Qut9�{̝�#� Y���r��q}�V����� q�n��6f������O������e�� �b����`���g��8t��A�ש�x)n%�W�7'��C]$�3�������M�s���-|��f��9��A4K�l��@F���D�����,��ߜA��[/"*����%�="5=�He;�^	1#F�,"�e���Zo�^?TV����_��z�^ЦE>@�
>�$�RtF��1~vu>'��s��K��Wk�pϚq���A?\7�~ϟ�_�G!
����&h4�[���

d�.����g+�񿩧z�N �C+�ޛoxt��mS�j�����;�'���kpڜ�L�]��)V3�� ���R"�@(����l��t�O�;���;�
Yͣ>*'�a^9&۫]�g�7p�v��W�&�C����C�ޮ�����lloP�H�l���(�����X����}�`���cZ��S���h݋�e�9Am3�P�<(�L��ho�|�h.Ϲ�о'C���F�"�ʉ苃��7�Jpk�xsJ�3I�U�X��V�D���6 �OfQ)R�R������r�l�i��Q�u�)��-�a�5���D{j�b���5{f����컈@����㠸.;����}l���p~�;(�:�6���,�y��{?%�9민
�8=*��I�)is��c{�{�#diۥ��,��lhq���W�!��a s��[q������%�U�?J(e(�T�sZ�%�����>��RnӺ��j�ܿPs�>��l��n�wEl1�u��O�!D�	B��Z���bC�~�3Px0{�#�PR�_�L^��,����A�ǁG�	�?S�א+}�PK   SH�X6e�b�  �  /   images/c0cd0a79-4e96-4647-8bb3-400a2b193618.png�YePЦ=�8����<Z���n$D���H�n��n��n	ii%�������ogvwf��g��_;��j
�x4xhhh��Y���wp�Ÿx|�	�a����������h�+R���k;Y�{��Z�yyy��stp�0s�z��j�y"A��F�(+����7�R���4�����j�����0���Ā���K���%h+˻���#�����SH�L"��8:c��X�d��˦��~����F'O�絍׌��~W��z�7|��;����d�CD(�Gg����Ȅ����S`s[ �OME��%��!�HK�VP�'�M����<���fU�*6��(�1��LH����u>'��?A��3, K/56���'���W�er`	�<5�WåvR���,�Du�b%�\Β�Q"G�Ni�p~ⷄ/��0Z�a���3Q%�`>x9�e�1#�b-�X��,�Mp� /�ɝ��� K�C/�*����&�U���oґ�9�N�#\������;ɼw֠u�PO.�s�V�q�K��= O�}�)(IH(q77��En�3���&���Z����[��n�:�9��İ������XYܞإ.#S��(CR2��Z�V�BXp�Ll�#M]���a�
�-f�*�&�үN+6h2l��Vb��9�"�%��Iʿ8�}NFA��友_p�V$�n�-B=���į+�����"��>aH5ğ����i����V�:ܞMpi�/�%�������0�Bh�I�e�uv�8��y��.*M����p��v�Bf@ 4�۶��u�uR0�f�JQ� ��Ǵ����\fZ^�9���7���#ps�:�֮F��*�+���g�M��}��D,H�����Y������W��;����y���#4j�}����>���˶�Z��g�K��h���Rǝ�}��dp~	�Z���=�)f�9��F-�g>iCb�4&!������&�ֽ2�����v�
��&)��l���&�(�	����ƯVjzo��2���{�����)Q�z����e�GU�����nS�US����6y�j�h������#k�EY�AE:r#��N������&h�U���q-�^⑼���ԛ����ԅ��I����~(���Q�T� e��0��Y�5�V�1�B�F�mo..ݍ����#;���>*��Td�rb�}鯻|��~J�擕�,��\U�P"^N������wT߶
�����R@�����9�b��u�pޓj+�|}�=����W/d��n��2os.�E
�k=+Z��#dK��)��m�L��<�a��gI���*^�"��R<��':�`���U����/B���տxNsW���U�N>�x˒�7��I8T�\#��5Q��p�g�4�~β|}������+�n� L��΅�?^CV��r�q*���6�Ⱥ_r��4��ѫ]�jIV�9������B}�((�������w;Z�ƋJF8��M�S[�Z�b��������,����Ju��=�a��,���ŬD���^-[�9�[�u��]�ҏ⫃�"���G��er1��&e��.,xí9�z
q��h�ɰ�i<�G ��0����t�/w"m?`M�,�m+����T*J�]N��_��fw�^{u��|o>vO#���j��Lg8���d2�&�Z��b�؍0V���f4 �~�h/ͤ��
_�{� ��A�I�9y�����B�K��L���<b��o����^ZEC���`�a���?X�5צ����b��K>�3&�.�
k��C�K�=��Pּ̑��j��a�RqF.�ZFЖ�-�ΦnZ��v��*zy�ag/b���@z(����l(����L�R�E�8�7Ȗ��f�0�9�nk\����5=^�����>uG_���?y<nP�@5�9����jw��>���a�6�Z$�?2�ß0��u�qB����;��x�$�8��.�sFy#��Z�C�z��R�
��m�#B�C���/�p�!� �p��c��kbdl^Ϭ�'�h�u����@w��G��q,�r���5��6,5R�w��������!A���Irܯc��A�_��y��n���1+�2��"�C��Pb݀#m���`�|�Hf�����F M�c�7vQ���ݏ�I/"C��Qc�3v:�J��:���j����B G?L{�hP�S�9,�oc
����w�B��/3�������J�ˉ���l&W\`�={�'
���]Mc���H�Z���p�OI�F�ۇ�[2�)��u
���&D��x#l����Gq�!*)/�*�qK�I��*lq��^��{数s*G�MRϿ�?4���(���@rs�s��]l���f�Xy��c�R�F�������SiC�f#�?2ښiZ [�,�9+�$jw��i������LV�	ܜ��'E�
�v�!"��o��}*<�Z>Z���0�l���2#	O�E�}H��d��
ta}�����	�����p��j8�����έ�8�4��'"��Ӷ#'�zT�!xY�6N�,n�1^PL��]���}��\�����1��)����m[�T��N[3 f'�2��[��:��S!���`%ۢ����"���"b؄�����"��=�N�BC��@�%A5C�:�����n�Z{�qM���?�2�Q/:j,|�w�f�6�.�-�f����l���:Sh���E���K�fg%�A��y�^ǔN�e�������U�k~��0�9�1�x�\pѤ�y/�Q�\2M�yrn��X�!�xG$=��hm/�`^V���Оq�w}��#Ǘ�M
Q�.���u�+]>��GQW"����SӐ/�!)b�|�n�ʹ���^�T�D�@��s�D;�sN��L ��s������hHA����r�N�u"VN ��9$����O�����x=l�f�X�I�8fWē�[�|�����Q��V�bl��%�`��������Y�&��4aon�*�՟|F�Q}�~L�o+���_R�#��'Ҹ&��-�#���L���'�����fW��ķ�!G�4bK�8Y-D~z]�v ����Y�ˆ�;�=^�װ�����<��n{�)n����BI�)���ltm�{���&'&|kӛ|�~1��3g<�
Aʈ%afs����$$xHl7��|:R������FY�6Qu��)���ӡ죢l>:��*4��?�bXcF�86ԏq_Q��J�KZݍs_Yg�_\��N�.����\�;�����-)���Wn��M��lgӠDjVT.�痏RěA��mk=�������T��>��oE�U'�6�ȖCLn�Jy�辶� ���� 	ө��a�[�[��?.�=�s�mp#��~�n��io���٣���m8�9Ɇ�GMD���79
&�ۢ���,0!Gl�ݝ^3ɕ'h�����]�����'x�
,�Uܕ7ě�w�wr�!�ڌ����z{q�\^X��Y�E��ދ;��[�p!m�����}�9��ˈ�6D�7��E��_����A��.M�p~�ap�~$�S̲���2W�}�7�X<6v5k��w6g�&����/��H��leIHzj)�Lt�fr�ۙ�ͭ#�+�o��������kԏ_����k��S���I�� �lVл~�>��Ͼ�]��疽�/��m�x��7=������>�-�dB8F��*�]� G������șUIT�1c��'>���������f4�fq9	��s�ҿ��d݂�)���]y�ELf:���(���tP�����gn8�}}S_u�JϘr��|�=\�P���r�oRE�Mo�pmm��<f��L��'�g;� _QSc�v���TFbX��G���ݾ���3[��w
���V�����j}"5�d��`9�x�&���Ϫ҂�j�i�S��_S� �g��b#.����!����Dy�9�rnyԶOZ�����;K,gR�2�T7�,���o���RHQd;���%��l`��z���vZ�ɴ�J>��#J�*�v)s5�[��o7P��
uޮƺ�f�pk	��{��;�Q�TR���(@������ę�w<���њO�o0-ȁp��÷���$��Φ��0�J(���ګ��z��/9�nD�_�j`:� �b�j��3h>y�5E�D��2Me7�.��np��ޱK���I�u��{[5)����J��}��O��-b������&C�I	���%�)��jן�\o4�1<Rj= ������z����K�L���uH믒�"�^�g� S.�T� 1|V����!LPv�!��$[ 	�������Tsy��WKvJ<�aXv#�I�t�H���`F�[Qz��E�n��`�L���m��PN�AAQ>�"���`Ѳ���36��ˏ>���f��d}j@�D'{�/h<�c}��s>�q�/�6�Q�:_�����df_���������P�&�:4��g#�����zx�(�>ҥ�X�w|����|(�"���*���R�g̛�>J�B�Ok�oD!�mH,�/fW:X�^g/!���]w��-wT���Jn�}Ja��2�~�f<����:����,�F�w����c�-�Ѩ;���*���s�ڴWf�zC�!�oQ~9��(����Wc�>�9Ue��T�%l
���M� +�R/��f���#��|oÈ����@��w:%FEi9�=�u���c�ceh�����g�9�������F5�p ��5ony��Ċ�ƑX� �I?��Y��<�M��O����˺OO|���N�9a�-�q�0��Q�ͦ�+[�k���1�����i������=۪m��M{)͵�uV�7Ƌd
�*8�hF%p�!�Y����V���Y9�)�����7���]��ޛ�ݮ0�"�0�΅p�z�R��l��+�Y�>����3W�D�����Q#�Z��e��i�05�Ԛ�ì9�� �R��������{1iR�8�wy�'�'��8�
�DX���A4_M�;�S�h��QY��}�e�#��-�m�X�!�V۶
��1�M���*Hj;�D������KB�O��S8i?%߼��MRZ��m�E�q�`ʣ\m�K�#>?v�[�Ռg-E�{f|%w9�8Fu�ű�����K�� ���c�����J�xhM]�e�:F��G�1HL>o���c6���e���a�{��aKL���鹲�Ap��8eo�� �������]-���Td 8o�{��M���q�c������-�p Xp�Lp���~&��ʭ�Q:psk�����c�Ui�/c��$KQ`�x�B���ϟ��?�:�8���܍��>����<��� ��$�Ga��D��O+������WSD�,��lCNP���6�7�ȏv���L��P����gxE&%���������S0zS�)k�%em3�
���M3�z��[�ī3�r���{l��1���hp��ՙ��d:���j7����9-�C�"�Χd���eߣ�z�If&0�\�/>c�BW��|P�x�Y�[(ɕ��H^�?���	�M'�������7?%ݽ�j�3-iW7}wX�z�.KP��{@�t�[�QC��I����,d�<r��i�7^Hkɹ�>0ا��ȫs_&*�~�ZQ���־�����=>�z����*w "r/`�=_��?�}��l]�R{i�x;Q����4J�Z���3\�����jh(!����K���x��
I������\޼� 0��+���	t�$�#?BzF`��3p݀��o2TT���$pKt�&�a�
g]�-W$.�����Yv��G�����������0������|d�qS�E4╬�3⓱6�ڒ�=���:j0~�l�O-m�C����ҺQ��*VZ��n�'�FQ{���\ld�B�ȱ��Q�:��+KT~�*����?�w��lN�:�c�Dh��Y����y�J����,$���Ǔ}`�~�������C;찤Ƕ�#�l#��&
�{����k���%��N"���}cf�df.�,�K��#�>�g`Fv4�O��9��x�9����?�6�?0o=;R��L@�����������?=�Q�a�k���fF����3GТ�r_�������@��:�u'��"��+?ʳb��x�'������#����C�a����e������}p����$���͍��&N���v���s�;H����$(��贒!�������FŬ����`V	l�K�5V��� 4X�G.~'�:��H,�9�&{�5��L$U��m���3M���빮�;��I��y���I���[}��1���;@���#Z�
���b�@�8��J{��=.�Ѣb�.G�+���_HiIܸ9�fqe�O�ߣr'qx�0)�p5�ʒD���¹�Ⰹë�Oqp��c�U3��Re�F..���ߐ��k��/�0	V�Jּ�l��~i<\��̼E�paTT`�L���W�
 ߞ��YK�_K�Ǣq�S���SI��a�\�,t"������e�ƪ�jGTNG`����˫�7B�Γgh��\'F&�^�/�D��˽��%5+�GE�B5tM�'���a�GXh'��s����՚(pFZ�I����e��0m�������?7���M�⛿���;#cU���[E�z���D9#t�1>��;�o[]�=�Rн�G��02�3P�`Dh�v��f=�Nl�:�^g2�������:�:������S`���g*w>I�%_����3`��RO���*�cl~���ơ��}إ��閍N�eg{J��N��Q_3~3�[��`���8���@i�";��h�q�Oov�:�_i���m͉C�k%�w��ǹ�&J���]W��k��b|��#� ���ny�� H��];.�
	��;|�}�eڽ��vV$�&������H��UĮ��c��8ꡌ�ߥ��GZ|� �*ז�N�)*�j�"'�DI��!t��/��Ƽl1�#��j�(��ي�ǧ��iY0]|I��C�#���}������;?b�(���r��̊��~(M����G����W�Ȉ��N�2�?��e:u���9H���E�u�ƲGO�_�1NV]��^$P	�7�[y J�Fb�(Z��Gh���� �d�W���-��A�Z�Їe��G�>��Vϰ����C��h�^��1q�%փq�5񣅨�����a A�9�jl��tflR���b����+9I�3� 	�$_�b�2ػ����M��Ӊ����wK�i<��7�~��yɜKR�G�1| 6�P��ҪotF��TPS��P�ӌ��C	!��i����D�X��y��>��M��ߋ�h�U"�,z���򭁏&�=U������.�2���AW�Ԗ�g�՘����<5w��i�\��H���6����?�?S�S������PK   SH�X~��a� ٮ /   images/dc707dc6-8489-41bb-a5bc-77a0670f90d6.png\\\S�� Áh���P%�lٲ�LX��,��
BX�Q���%�A@�� �0Leʎ�gb!��b�����p�=��y�sB��#=�=�{ /��E���-��|��@�W�]~�a�<����7x��粅"������	��Q�K��&�����N
%�����p��I���%e^S����iP��`ȓ��P�ej�l�{�y�o�!O!rݢY��بߚ愳����}���r�Wk괡XY?�q�?�üh���!͵�/V��xt�e~fc��	�O��D�:���s��;%!�E.�o���˘��P\hV��rɘ �;����TS��{k����EA�n�Z��2���|��k$8V�p�N���$&��������Q�9�HO�	��T�{���M�*��o��f���̑��M�<�!�f(nQ����P/ h�fvh̜�,`�*�Kp��e�Wc=W*&���s#�pSx���]jr������Y�]`7�핮��jʿ#˰?!!�\Y0jn��D� ���Ȳ���h��87Mr�q|h㡴@~�K���g
�	��Xy6\���J��ځ�ӏ�u#H�u!�}��K�����%%%v�ou�V'���'���$�
����vv:o��Dz����p��r��gD�*������Tc����u&�17Jw-16������p%�8Ec��Nl�B�{Eُ��^�LG4� �s3�Y&Gބ0�F�٨����?l�HIƾ�䦚 Y��q
؜$ȁ�,S���fDz|�e,�q��傆��Vn����@>$2�r$t-�Q����a��o!KʐĦ���H9�mb�����m�Ž�u_���is��=ۚ����1�r�|ϐ�B-a9~X
j�MD��+	��#ҍ�֘	��1//�����")�	p[�e�5���(ۯ�N3�� d�)T�����ɂ:�x�f�h/G���%�����	L�e���fx{���}~~~��J�1Ε6/c�&�
?LDD�˓��3�{����g?�eB���Qsn>��>�2�+Ȯ�\\�1%^�+���q��>�n���R6��]�]z�}B�u\����uv�Y��H/$�W3�
&d��Z��v���#����ї����k̉�����ڱGw4ʂ��W/��� Ɖ��OP��m�*�E"7f�TU�����a�@���+���=�o�a5sTL̖=),�Ek�k�:V�[o�_�#� �zbўׯ�o��Z�Wud��x��CU/��Z��,L�s�ŉ�kY�����"NN�9�s?���ma�����i�-g�1����H$_g���d#0[��n�����S�Y� ���>snBj���ݗqt2�0�׏�΁J�����7Z�|�2��_���R�t��� p��Sй9;��q`;6����@��VhS���[�0��o��V�e�_|B���l\�Qq���So��D�����[�m�~��B��D,|x*.F�Ƭ_�8��J$�Asp�y�f
<�]U6��Ka����n�����#	,�~��=w'H�g`��w�z�<s��@���Y�Y��F���#����e^w ^*����&���'�
o��$5�8����j�����	^�,-�%z�h���K`�kʋ��Z��**����J`�W	����5��#��i���h!����6Q�#l\Q�¾��%I�>}����t�=y�y��~pyĒ;�H�Xc�u���޽{ͨv! C'����|SE��u@��;�u6.^��~pG��
� �ژ�m�@[�:�������EEE����G������b?�*���������6��7)%�iv֣j�kP~�Ӑ.�Ă���:�tD�B|{B�B��Ǭ�A���*�m^Y	R���_
�~�VP@���1���(g���l����ˤ�E��m6����@��:9߹���п�YL	�i:��fdZ�c�Z-Eջuee�KY]���mUCEUUF�VT����206.���J޲DvM�d�|�v�3l/��i���9����ϴ��Yy���3�;ǲ���9����vnHa��zC���d�?�{w~��|2����r��,D@���ͫ�P�[�kᅠ�,1z3��@Sd��o�<��Z�x��Ey��(韤�����H@n��̮��0���k���TM����PSc���q�h��m(�Y�
-!��a�؄c�o{�����;Ϫ lv�R�
�eXR9N��6��c�ݽ�j�y묬,�/����bF�a���؉����7��Bl=h����>�n��P�J$�\@���P�y�m����_g.$%'7JTc�e�NLִ����������=�g�'?6�L��U��N��=��g�j4B�- %�O��@%���7U+D���oM�"\�"$�p�� {��+#1���G��P������G�8�f^U� �!߆P��ɲ=�Lb�ض�>6ʎ5��-�m��X�7�E��EvQ�K����(�����- E��ռ�*���к�01>�s��� ')���.Nb��̔�98�p@��b���w�X ~*lD���w��-����B�@�=v,Wc��=�M//Y�o�+����R�U���^_�&�}0sD6�h�I#ql]E"k�뾤�bS�4�]��IU�l[�I��^�7���z�5M�뱂��@��l�wTh���8�4i=8�j|�ߛ�8I��
��$�
�}�{<ڄ�o7�C�+S�$�qU#�3�FFF�����r��ၞ�Wz1��c�N�M�cQ����}�".��O����*m��A_��o
GϚ х�ie	+��dH����Q�kE=$��m�2�0E��趖�`;���8�31J���̧(3�ۅ���w���J/�:��K�\��"��PGe�m��=,����Cj!��W�cVXU��L||*�'d@��������Z�2_9�^uj�B�.+��!1���RݡY����)�&)>�B�פ��HkU��k`"�c�/�oS"���ʦ��6C,��x`����vb^�p�`�Q�Ǔ\lsDY�x�,P/}��r�-i���Y���5dx�w8���t���6�#�q�n:��������f�de��=�����Ĥ6)3=A��\&�x(�EE�f�z�����FWG�l�2�����0�㥒���E�i�^��QV^*S� B��Uqк����P�zK�'T��I|���	Tb�&��S����<��51��W�H$5��(�>nV��*
x�Nh��@�/DDD�$n�'5!����<y`3����l/`���O-P�>��-4�һ�e�U|�\�
�-<idd���v�Çw�����<��[��Fj�f��������L��Ӭ�\�:a���E��)hȵ��Չa���J-���`�[0,�)����
\[��&�,5U�����JT��;6�6	)���/�^�� ��gz�s������]��`w
Q���J�����>abA��V���rkʳg�)��:�����wL�^����6�� TT��B�b���9p٫u��ۭl���2��C�uX���_#	���ڴ������c0�N�����{�����J�H�(�aԏ�Ƥ[����ϧ� T���n.I������;�F)rh���bi�
�Cܝ�޽ks��qF�G��W��9�o/�W�Rm�F������'�m�(&�M�h��z�4�0��z�n�<A���(o���]��4����a�<�$@�V ��om���Ź����+X��H��ޜ��P���~P#ʸe 7�v/��k�4Tj��gߝ���8D>a.�`aiY58ƌoP��UO3���f�ח��/K�j�n*�{�� �@Bv��πn����w-9�E�mL����S��0��/.���WN��_��H�&X����Hnz:�:;CσT�����ׯ_����ۧ��V����K�G�۹��K��>-���f懧o�v5�h>@��'3�a������f�ֽk�mv�G<�S>s�С�xĪ���J�Z��M��k𙅅�)����6 s���1K�^��@�z��ʵ�*�P������"7�rͽ����S���q͹!5`*�/Nu�n8�+��4`�0>֤?<������[+�/�?^\{�9�F㾲�N�R�������d��Ҳq}-kS���sֶ&t�ߟ���N rMJM��Q(:]|��}J[��r+�G�	]�E��]\�JlJ����5��2���o+���T���|�j�R��F�Q����v�\x���%cn&�'l�nP܉��X��М`��C�����Mq�ي�@hz�`�KЪ�,��Y�{�III�2̭mlFD����g�*,�3�=3�X�ؠ��i�y��0I�����P�0�v��qUI��.zn�p�f ��a㬉h59�f�~�P�`(�	��D������,J�`Y��G���T �a���c�7NY�{��S�;�e����3lgL� �s{N�>����$�5NN�Y�%@X��E��A�L�`��``` }����?}��xWt,		��8�
`;��	,���NM��W�^��	�`��v_[��xK���Z�
Y����W���eƒ�@�;���+X�\��XfyTX���C�꼩�o�gwk��oS��I�/����ơo��Y��Ü"1�<�"Q���_�|^�����TSZf{K���kEӌ�'�2j-o����������n�9��ھ��(M=�%#T�c��
V��%�!0ܲ�ܜn�*�ӛ�|�`Y��� ֓�Y�?��-S	�t�&r�K11R�Q֊ ���V )P�L`�����tn�O�֏�#K��bmY���Wy��`�:��#֌mpE銰ʗ��1�!'+�i���>��Y��tT���@�`"k[��%�2����0�nG��L \X�x5���u��4�3 V��`h[�V�L�ri�{K�Q~�E�1\�7�LykMU��+ �Z0��tʷg\Ē�ءj}	DrL�45SY��]�i������B�,B5x�s|�����5�!	����jz���?���m������	�X���2�JF�Vh��>���`靵�_X]��f%��}vu��o $�}���6��r5q /,�Fy��N���<a�
���xS�K��4  \�C5��r��/7|f�}�U���ɞz���Z���Y[�]_�ե ��߿GIlMȌ�p@〩L_�0��r��џ<M��}ZV��5RO8�t��.�@�w&E�_X�Z�T�,,\[����@�W���M@稠`Uy���7����h�b�S?��G��B9����~�e7��@�)���������]s��a��Z�u�z�$�{��$3$�����COh����ۦ���i#p���&J�!�;�\���f?i������E��M�gj��7�OH��d�rйN �`?�Z��x�%)[;�n`����O7=����޵��Ngg��_6���~�rq��'&ZӚ@S�N~|�8&�v�'��c]��K�W��1��4r�	�\<7��Z���߯�>��X���IFݯ�mۿ�l�.k;���!	� }	��3�zr�{��]�"p���2X]3����5�N���K��-��ɩ�[k`�Nͬ2�PXo*���r�y��P��M�A�Sk@��=d���*�D.��'{�Hl,��A�� *��.=�zs0̑�e�oQaO2@���U��o�,� N�wG��Q�'V_{s̰�Ƀ���6�⥒ң��������6�@ث����#|pI�e�(��	8k_�g���C-tտ6<�'�W_�p�ڡ���YAM��&�jSب��}�_J烜��X���l���S�n�%� bSk�P�1ߟ �he��X����<��7? ա�8��J���X����k��<^㲭i"��۱���S�A�M�T#rrr�D ?ы�\g~�(QQ�fV��O%���,6腟g��K`��<���s90���4X?�B=����/,���~�2y�a�[�� /Wל���!UY6y~ڴ���4$�J������u�g���W�}�8Q;^rݹ���%ǟoO�z���U�}�:[$�p���y쓣<��bmi ��������?�m�-O+�T�X�������u�2�xs`p?@�C �c��B�R�m`��0<ˏs,O�V�x�$�C����c�'V��[S-��K3�k?>�Q#ǧh��8~qnC6�������\K2�L�h��X��ꇶ�˓�C��Z�ִ-��@�Z�E�Y�v�5��1�ָ+��-��ָ����%��E�s��&��s/��� �mqwb�X�����|a�~ds�g{�B�DA{Q�Sqc������D�]���Z��,�)��y�X�O�-��<�շ$׏�i5��ʡ`,\�87�Z���n��`j�\�N��.��o���E�����{�ID�$6��!�?/"6{���a0Y�*�v��_:��ء���~�.��۠f��a�c���B5�:��ڶd� m��V�d������/��R�й	�����/P[uC걣���\Ǣ�H6�e�ϫ�J�PuףF�(#Fk�l��� ca��/x�����&�=��r���3�!uQ���{����J�>Q�ġz�h���I_+�1�L���C
�A�h��C��\m�&�O�j��P'�uE��)��a���������˾�ޡ��r��SbƢQ2�1S��ݐs�;n��D�m�Nw2G�Y�!ayO�O����dY,C~U��!z[��K�����p�<ۋ�|ܯ+��0�gϨ��m�az�	���5�{�RMY� �$�lz`tr0�f�� �G�v�V����:�_���Ƚ]�wC
������r��T^n�Q'���n-�xM�$�����q>!^�h9Q��c�@nא
�Ճl�n�_D�/�����g�k�a�2b��b\�4� �?�e�N맃E�D+����0�j3F��
vz�A*_���p�\�y�;o2nt��.x�9�qAa���}�1��J��
u����$��&ɾ?q�h���}Mؔ���2�����۬$j�_�[��A(�;,��+��I�7��A�Y��m���++�O��,�$�d�����ȡUFH��(�S��:U���w������!0��FͻL�5�=�g��vx^_�Jv���>e�b��Lg�V<=_�8��h��>y�0���61���j�O_��������@�X�p�:I�2�qm�/�}��RT`z7���[�a��V�bSL6��ˆҷ8��7�WUH�]t�PI��)c�1ùw}`��[��9j�:@����1h����[3d�����{"4c2/n�j��;�aw�L,a�p�`����y��C��c�kT$y��3�����8�:jR��e�	��g����`t9
׵=T��
H�w⨟(3֧��������Ĵ�1�Q&�m������߁sHw�7��1�	mK�m^����Z��rA�y��+H�b��j,NO�n�"Į�HJ����s�d��!}/��6�Š_@u��4 ��w��(μ�4��Ѻ�#*���t,0vRd�8ǗC7!�v��>�S7�ǤʑA\I�3?Y���H��U�y�&�v� ʴ�i[bp����;�E:��:Z#&��a�ua�W1ߒ��HUY����ˁb��D8�_��W��e�����eGL8_%���ȉ1�$oWu;B
�?�a��tT���Xm���ޮ��:K�pg�����$̺�w���!��vz<�:KΎE+��j����qj�}J;J8Y�r����B��t��:BS߼��?_�Jt�vMtGF,�*,C�p�G$]�	)���ȵH�͟�O����!KOz�ۤ�Wwzn_)W?(�OG��>-I{�N�)U:�a���;i�l�jw^�/�VCA�]��%�W�g ��/ӟB3��7`DsL�$9�U���er���4`փ1&��Q旗�<$�1�3��`.\e(��:��*���C���3��ѧ���"����N���=؍��%κ��
+R��8��čA�.���2�p8�Zo��tO�v�h. =X��	;�^X������`��G��v�����e�3&F@1���`�������A��;D��0m$�0������/�z�}��&���60յ�� o�v�O�*%�A��ݳ�bz��K�v^a#e2h�8j�O��`+��9�v����O�&� ���T� oA��&G 7;����ϒ�H���ə�Ab_@̏�h����J���/�R 4lg>����Xкщ���̋0KV���.�b�����OF/z��B�]��#v^��1�3�8N�N���i^������xЭ2��dE�+�v����@ƨ�(����H����L>����g9W�1�=��i�Ϯ��o�-M2��L�+uw�6bGj�� ���g!�۽���N�����#��h���!Q�!��w:'�ea��Gb�YP<���W���<���j'���@��c\��uŚ_ND(_�y�[&�O�b֯��p�9���-���´�1�7`�]'x"Rv"P�N(,�d�%��,9 ����(G �XM3�\�����H�;X���Z�ť����>l�W���y���?+͇^��)χ��?y�9}e�yZ�X��$��c�i� �S��Mi�}6~�A�)�����qh����!I)���	�1���9,L�<lL�@"��8�~Q� )vdd�*��2k�Aɀ�p��H��SG�����!���p�M�1��Q,SHCl�P��x��^�tG��_�6��5Ka�b��`� d���/���y�L
,P���0X��N�K�bg�u�B��Ǝ��D�������G�Mc+݅����8#�o�&�25D������jV~b�u�3?y��������$kY��y(��G�01����u���hA�0~l�����ql�ߤMݑ9��2$"�s�h�]N?���D���Z�#��������D��k�:�8j�yۏm��([y�d������]��z�����ioxԐ��D�6/aj�Dk�� �_f�/SFM���l��s	�ߐ�C	�C��v����V���2��5��S�|�����XX5tNGŮ��SE �O[mC5=����	1�n�G&�ô�{���WN� ����'$���o)?�QXH82y���g_k��+��vG�������߂{�=-/���fk<>�d�Obnn!_}����o��r���-�rl�����d��p[O
���kz�����P�W�/\�-�=~��4r�=��_������?�|y�TJb.��H�p�)k�z���i� �=Pأ�l�f�����(ͷ��)p�?j���{��۰<�j����ϡ��צ�g0������\��
� �|��a�b0��\�;,ƕ��8�s��'7��szr�ߞ�M6��>*�6� B��<��9i�N�}��u�	�%�ﮦ���%Cs���$�Qҧ��jm(&Ց�L٩fl=l���8��;ҾlMi����W�M���E+�zp���� �?2��摕2�����[-�Ӯ�_����B�{���W]}����E�H��e{���k��>5]�i�W*>��H�P��ݭ�G)TD>c��R*�����#�ɐ�~A�Wr�͸�x�_t���T4�/�׈v�����Ԁ)7�Lo唏8-"?Xͩ����o���k�w�'�y$2�����,�����Z�b�ٌ%ņ:��s�N�g�)Ƒ����(1�M��ɘ���Z�q�q�EA��{�a�}Y��S>�+}ͷTB�(��T��"�&�Ά��}6��>�}�;�JH}�[{�(�ϣ���%���[��!v�j��(��Y��__t?��;Xȱ"wp�+���3����kֶ0Bm�0����1���q2���@�����I��g3�"�^�NTŝ��������0ب���U�0D���7���aK�F�罹����g�+5j^��q=|;G�= -{�BY"͜B�ή%�,����^��o�l��I��HF2��-1˭�]����=�o����}D}7�����a�߹D0�WЍ�0ą��%F�9�2�$�ך�:h|%�y2������rYHJ����ڌ�)�鄲�|)c�쳻6�8'p!q[V׃=E�;L��K�Hi����Y�G���:��[^G#Z!)���Z�@8lE �^��r��ݼ�C��4}U@#H��*���Щ���W �"H���v+`�T"���/�3���8H D���p���ri�-h����A�� ��4<�X���k�0���u��A�]�<>J�����3ag'2��� �����V>����߯��m�&)�Q�H��r�L��� �g��;=�РS,S^��8Sg�u�G&B
 ��o�d[^�=�+�[z =��{���e�ο�Wj��fa%�>���ɴ��ڜ��i�*zC���Þ�x���Y�o�75&����];�:�
�ŵ.MS<�ͻ��5Lh��M�vi>N��ﲽ J��O�+[�¢θ�*�7�z���yv�%��a����Ӝ�P��Ϻؔ5����~��MDɽ!� ��0����~li���u	Z�AmȀ�sV_���q^���O����N��J3���#��m�؊2�!���FA�n>��N���df�)|z�<�>>��$��"rO���M%���&s���32�1�=Ј�����Os׿���v�ushD4�x<����H����:������-m�S-/M�/I�
�szq���f�@�M��X���bczg^C�:��/�����ʮ�]�f��0����U�	vmCѼU���D�U�� �v�2~��O�ē��ǡ��.���(銎�����hкL�_�U�်�G����^Q�O��(�pT�����]rf�	��Y�)CG���\�MON�&��U�Q=��ݯ_�C���>�.�p5)=�98X}N�󮺺z��R�vF�nC���U�lՀk��I��p�u7�u� ���FS_V�!Ô��so>==ݰ�Z��9��E����b�F��<�%���Q�W�W���f֝NlRް�E��.��ux����o�ᝨ�E-���o8-� ���t"~?���jDJ�D�qU����'������+���#0�3ٜ��zz޼'ѯ�|_�H��uN�������T���kB�(�PiӕCU��3)_ߺ��^��93���X����ٳ˞�����4�k�}����!ct�����1]�/6�a)��R��~�ʸw`��x���'/���.�����xe�n�miӓ�'999Y�$����7�/!6������N��8� !��̤�%�u�����y^�6��YNWE� v������jЎS8���dwGxCPl�Ӿ�˖����̳�u��8�3�[y��Ŵ�͛|��G�$��W�X��,�����ҥc�G�ʌѱ$F��F��,���ʙx�!36�D��gm>�t>���~��bFb)Ԇ}�kY����H +K�ԇ?���@%�@������D����-h��E�>��psE���"1ؒ��v+�����	�,�_`��/М!��h[5W�=x~��	�Oќ$��l�9�:"�Exl\���^���kV���o��l��:���y��8�G搯���3�9� U>W�٘�'#�>/>I��2��{>T��I��!�aBV�c�}��|�PݯIG�Q�Hk��Ʃx���=����h��������Q޷N�m�i�}���~��Ec5��ƍ��"R�?�˶����uO5�@li�4��oyL�Dʦ�vJK����9nF�[��{e)ڕ��������Y��3q]ۺN���͹�WD��
����X��̺W����լ�
�{�����+����3�cqM�b�q�[�o�}B��Ç�}N�&b�����7�Ż��8�+J@+��g�� l�s<�}y�=�Ϸf*�;:�<1�~?�*�)��$��,��(l��P=6�<n�kk��<	.
G}+�=�Μa}L�]���ށd1�!��n�>̪�s���>o��2h$MD���Dj�׾)	�k��o��?)�$Bd-�?ݢWg@b.�t�|�!:�t�	t*��L��s���Q��$f�79��&B��$&�4�6*�uZp*^`�M��)��aa�	�Esqǟ���β�J�vp�T!o��#�'h!����ğ�$��]���М��"?��-��k9`���q�����BeG�K+_(��8�����cxY>��1�O���Op ٘�W�b�PS���Vz����U�oj��uU�.�c4���sw{.ތN	��m$]����r�~�z�L����|�uM�e��u*��<O������L��11�H�3A�mUcz���HʎH����co��m�8�3��.�>{i��/�p���7��Կ�DL]�EtP]]$i���Pl`ĂA�u�����ԗOE\OJ\r�nN�byZB����\����Z��CS��sKh��9l���3�^jn�?�\���,#�Dz�#��Z`�'nPBI�S�K�'dRo�l��j`I-X�j�7�3>�[_ooR�n"ayI~.�%�����RNhe�3$@`�O�k�Z4/r gyt%Dr�Wf���׻(�,�VMryqE�&�}�{(����	����' B��^\��{8YH�[�$_Hf�{?��c�R�kL������0�F'��s������NIF���\{�����<�˖}�s��U��)W�<-��#��&@�$G(��܍��DP�B[��<��@J]{��T�B����ڢ�#83�镴U�tٷ��"ü�h�ZyCv=fӈ�5M���hő�ˋ���mӋ���/:uޓ+"2��PP6[ͅc[8�e�����>�~�������δ>>ӢEP2��|�7�w�k�
�}ө�y�p,���S�<����R��ܛj������w��_�T�B6�tH鷿[�XEx_\yų%UN��]� guv�_���4C��φ��o��Lm��U�)�@�D��d+x%������b��"@�lv�����IR�;d��!���^�����In�B��4i��S�6w3���x#����U�OTG0�Wწ��;88H�U.(U��k��搸�Ǟ�����l���k��sY؄@�1�*�J�R��^�"�/���2��:����5��p؇�M;(kH�������d^���/b0ݙs?Z<�Ry- ���������Ч�����Qw��Q���ޙV����I5$������+�%g�S�b���n��~�qe�(淞�*�ȗ,��!;R�ҿێȕHl206�XX 8Q���1��c�T5nӡ���ȦR�*��SӔj����:0����hI��2$K��$�N���>t��)��Sq����۷��={��u�q�)��~��%������=1��)�I��xS� G�-�?��pN��Ԗ�����4���,
��-�r�1=u�g���lC�}��E�u�ԃ�G7��i27��cҎ�{��Y���Q��&̚kW��ێ)�4]��E�{`Z=ǖ�{�7�NI��X2�·��D��t<H����%v�~�^�����S������ �X�v!4�T����c�#���4�-c�j��3�ʗ�bO֯<.��dT�DW�h�ة2��Ə
g�����=|��|�����l��|Y111A���n{�B�ȱc����Wz1b��j&��"H������,մ��`���Q���6B
�t���Kk;K#'9x}�Ћ�/�M�t��/��I�N	��xC&�Aȼ䪲��zZ��Vr��7����u�h��n����(������G���z=ο8geulnn��W]�>���422b`d���+27�,��I�5�-��8��[��K�8z�͹�-Ȱ��+�w�mS��l>ϣ*G]���-LNM��l�����L��Ż�����}�J�Q�n���:�d8j(�C�c��P����-��-=�% ���<YAJ�t7�݇V|��V{���߄)=�5 ���[8���|����]��G��Y���@���'�kJ��텅���r�t�(��[�| �
��:}j=��e��$�;��g&ք�[��?*
Cph�UK�UK�j.㯜��b֎r�7���}!Dp��
�R6O7�M�k �b�Z��9���1�{1��	���@*gخ
Π���3�}�iڔ����h/ |`S�,�o��L(][v��;8�J.�e�ށ��1_;�1��f�F��6Θ#����&�氯^�����t\#�qQ�|�8���Z�.������R.?�vY,V�7M�d|��S�5�C�M2^cb0���Gu_����d�Ӈ��F"�bccn�K|���_��f�U�V%E4�M�� �"��$������6VI1���|w�Zk��`Ւ ��Ix�F�#�}���m竾wa\����ڃ޵�y�!���dn �-�ڴ����@��=�p��al�n�������O��R(NO����[���=
m,SM�>���ܯ���.Z׍��:<q)o$�8�PTW_m?2��j'�y:;;�}�c���7_(o�z}2gI��s��Z�ZK�|�"�|(�^:�to�+�LK�?��tlJ�)0*<�l�eڻ�y�Xd�35Y�J~Rc� ��~Z�U��(o4lA5���\��G��)��$cX
!�����W���z���͑�G�U�%e����[+�ؔ%�.�}��X������VO�-�N6Q$�=�0�Qݩ��乸��;������� ���@TҨPu]к%vU�e s�I�p?�7Y&�*%��fL8 �e�^�6�����o�2��=I�Mxw<�7&��{��8Bҕ���^4�����<���/F3�8[;i��t�8k��P���P�K�����-����ص�<׿V�;{��; ��y^�՛�Gss	�U��MdM0�{����u�|��<�;v>�=�Wy��,����oyY[�n1uݼ�v�Y��	`��uCa�:R e�t��X�M���\Ȗw1�&6���[�����|fT)�JV��z�6΅��̱���%_��\���s�Yw�$����sz�������;R�UKi{� ���4Dt'����� ;(���*# ������FMf��o�z�0=���wz���}x��`���w[�|��xOrƥ������0��5s��D�1���rϦ����8��zR�⍺=���~f���[��� 5Wx���Ytmk)A���wK>���V3W�O|f$L�XD[9�������{��l^uҋT�Ƚ�CH���k�B؈Ɂ��.A��L�>bhH�Xl��]��ݟyް��D��O�(�^�Y��~�]���c���֯��%��e ����{翼Ɉ�/FQm5����'�$�``���1�ɽ��|�,�t�@������9�\g���h[� ��d���3k�yJ��D�"N���u��$+ל�T���LF��I3	�Ћ2\\�{i-ۣ��9��7�	��-ة�����t�q�ri
]�"A�ȹ&�c���`���`胭#=��O���T�=���0����M��#:)dǰ[���#�V�T>a~�Ź�#��m�)�	�{-O�ݬl�!�0��R,�N���ʙ+��`��w;t��.[���ϯ�h*(���((�}rr2tI�*�@̯�����JG};�����>�M#\�s�p��m��7 �-}?��vgؽFtm���D�쒋�3��ߢ*�Gt�����g�}��_��lՃ�=��Z�.��}�ֆ+����ߏ��mgv����7F�\H�@���n�{-05�N���I<��D�q8�7چj��r���1�9tD�s@��@�����q��SXӧ�i�H?+�~�����T��������<�J�"sM�;Q�|��YY�#d��.`������9�����`m�*g��ܑ9�UZw}�>���][0ӽ�yW�J��ִZ�u�<jӘ�o�.I�n�y*#l�<�&�V����9�L������1���.������7j N[�S��@��myfw��J�G�@���EF#�3����w�ҋ\{��5�J)|��;��'����K5�W��4��: j������F��	�I�?�jP��I�3yb��i����=`����/�>� ����=N��`��=ϓ-�4�����g먬��43�8ywA�뵳o��C��g@��� ��5ꔼK����8��qV�����o߾������>D5t�����R�e�Z����3���kI�sW��Ԛ�m\S`�Oف�(���1qq�CFY;t?ۖh�-����	B6q�ޑ��˨�vZ����S�G�� 3�TVF,�r:�1Q�������]����O��X�,�,�o��aٮ�ȇ����V�5]^�1q���!2=��S�<�z��m��jz����>��~� �G�qh>�u���}�j8�q	��2Qb��x�����^�c	�f\�&���lPI~!)O��m�~lW�KL��� d����g���\�����Mw��Qr,z�j���5�X�QAAvʿi.u�H���+)��� (J��CL��h�摊��59���S�@��000������]�wo��^�=���<�0�4hF�U�IѶ��n�6-�?��8��W�_7���D"l>��z_���XZZ�q�gb�y������=�v�c�Ho�J)%��9��$�?~�/�XDƮ�X9}�	�]@����.�����xY����r-[�eB�d�ۍ_��+F��]N:q"���o������ֲz�a��?�����Mֲ���U%�M���t�*!H<���ag�  A���ޒSS�ǚ�Xᣇ�lu!�.��N�*$5OQ�J�V8>�es����v�j��< �E8/9LA��-��>V!��M�~��߻v�ĵ�$��rv�r��$ Odyy9hy#̗�/NF�������Ϯ|��t�3 J<"�f竾�	�a��+1 {��oY?�$��$�Ν/u|�����U����}��0�����׾���u);U�%�)*::L�~�ڞ�Jw�zj?��Xc��p����S��9oo9�ȰT�|��Zeo�����%�d�qL�B�w�b��sm=�:�a��JX�;ݞXz�3{#�Zs::: *|F?�>����8��7h�ug��Yڥ�#�p�ͫz��hh�=����-rh�:����wU.~qcmMp��8�E�D]�А���m�?Y��Xp��M@C�p/�cmPd��-;-�bd�Y��rH���+��[��R8d�g��YB��$[8[�&�~�2�xN��x��N�<�ԇ�C��{}y�, t��ݞ��"�HK���嘪�h�{��?R��>>O��U���LLL@n  ZsL����I�N���J`�VI��u|����ś�}��|��~��3y����4}w<������HV��Q�){o�P�̮d�ۑU$:V�)#d��1�DI����>N�ؿ�����q�sw�u����9����K��۷o+�c����jxԝ���^��j���mO7�*��&Db}	A� ��'���l����Ȯ��Ȇ�_�i��9��	��.�7��H��h���R��ǌY��b@��zM4��Rʬ�S�&:�:���)��qb��O��Ƀ��>�d�r���3_4~��
���J�j
�
�7b=$��ĥ^�: ��,R-�S�9�+]6�s�0}o�h���r���g��X�+�5D@"&���)���ʎ$�����4��G��z�w��"d_�~M�r�xH"Le*���Y��[���-�Ժ�x��Kz��ri���������{.�Ba�7R�⩣u<u6���7���ɸ��No��6��0�0�<�X��MZ>�a�(
��Ȋ��2������N����P̼;�c��a�o��/��HXy)y|s���=�d��	�VU�K��X��-xWX3i C	m��i$	PW��dI�CF�F@����Y	�}�F%���:Н�*���&�m����|-�~�a�g�B �=�2}}`���M�^����0Raa�=Ț�pl��WͭF�8�ח��lh���h�Z��R�؉dg��S��]}}u�)r���e�s������6�!�M�f��ք�T��X���0.@z�`����1���0v�ҵ�2���T����j˶����SW���"N��P���S��A�k��z������;��謽��e�)��
v��$��-^",nG��TK�Dw��8ϝ��M?L<���A@*i��=1f%��%r�]W��@Zk�G
�:���F>�=K�!�J,t�.SN���:��U-��#��/:�F�n_�񵛮'N�ɱ���V1�P�Y�iW�۩��_Қ86A�\.'�=xU! ��N����g\��I���T��:�:�ם��_�#� P�e%�`���A�?Ra�3�P�- h�4d��Fg�KS�y��^j�#19��=�R���8�d� ���{^�m_��3�$�c�|�zu��7���C�*wBBT�aůݰ�21XY=NV�\�L��%Aqpi�gV���'�n�"vK�����嵵��ű�z޿��4�W~�jjf�d�l��m��7�E|��0� m<<*l�h#�,�kkS������E��ݱ�P�nn������7�sQ�(��Z�ݥ�\�TV����Ѕ���((*���<j�a߲l�p3|
4�ň������=&��yyy_fY�9>����<<��9kSO�|i�%�����w�G�K_;��f�L)b���Z-������c"bq��e�Qܐ]�-�!����ֹ�L�α:�%k
�O�kg��K��XX@�O�\�=8hȚ7|�R�htՌ�H�)����w=}(�G�>�V�;A�����w����bꕦ�����K[A���s��!?ޤ��)Y-H�l/w)=F��B��k�����;=�cn����N@���
�̋_jkISk%�Y�ѹ���7Qi���:1���Η��T<?{E���U����٢��v����Dh� ��oݙ�+�T<�������BXbB<@#�LG�$
�|�yt��8��j?1�e|Z@��~����CK�Zh���t_jl���т���[5u=0 �����h�usVK˭1s�5g��x���c�����\�2�ՒH�������w������^��~���X�������TknPbecc�l#v�a��$��7���1�� A%����C<^���	X����\dGG��u=��M{��^�&_�yQ��y�e�`ޥ���qmZ_Ta��zp��2��{s���A=��Y����%���Ö�/NB󌽩�i�K�&�P�Y�3ƹ���4�C1�W�!2�ٚ�T�K-;��x�qq��x���Qw�4������hσT/��@�G�8rz#K���qo���o��A��8���{�v�LF�"�'����]Avtv�J���y����.��H���x���(٢�M%�[�F��E���$+5�΅��kK-h&��V|�����+�R_m�i�)Nω���(̉����>>�<0 ��ׁ��P�(_���rTn�9�J2�IDs1��'6A�N���iLqޫׯ����B��z֝���.��7@��݋���x-y<<�D�kg�Z�}UUb��	�k�����	8�V\H��OLgI5hb�L�Qw`�j���P0�6��c$��7[���Ν?��l�����-%6�8�I�a��	,'[��h���\����/r�ξY����^�SZ_���+�+�D�ٲ�$�K������3��:D���k���?���g{.M���z0&���rO_��$�A+�������)���h�1��0ڲ�G8�n�@����!CP�P( #��R�=��b���y\S9^�~�b�Y��߁&T'�|�G�,z�I�f��Y(��v-��������u��g�4�C���Z��r"��g� �W�V�N���Ъ:��gF�-�~�8��;����z���Jի�ݻv�͠�;���k��H�1��~�{
�p����h���[�-��tQ�w���R��?���vv��|�6Q,�ÿ�����D�7�:w�}��͸흢p�K 
��G�ݎc���4W�t�=���w�Q�P����
���X����ͯ��s8X��B��>�F�����jdC�eb�\]4�ąN��/��Y��`*�s���m�EqR�R��2��f�(4�U\���	P�����x��GQ�
E�m�]D�=��ڀؽ���'i�+��tޙ���ӌ�;��TKK}�����\��gJ��\ZhGy��mv��S�jyd Sd��C�~��!%������.V)��HJ��F�����<.H��z������7��s�^�*�G 9/D���lv<�.�龹�~w���=z���6���%=B����0ۅ��Ҏ��{@��j��慆Z�Ǯ����j�v
Vy׹�>'��5x�EZ�	k�����ޘ�{�T��9���K �G�L�՟RY�
�D4z*4X��xj�5(����7Co��Ih�JN�o��*�����_� ~�R=�e<,�,݃'v`�LB��9����,���-��M���qj ^�~�/������S����?y;J������=&�me�
+������s��k�4�j�f���=������T��t����??���.Pϼ��ԏsZ�b��=��T�՛pZ����*�>��j��܂H�FMo�/��I,j�B�D���"̓BִY���yd�ʛ!ĩ�9���C������cT����⧶8#&�r�P������ڰS�-Y\s�O5q����Ai��$���jn�0�bTl�����ϩ��v��+�nn��3z��/���r-�6ȸ���}�x����꡻�����nMMM�-k���U�<@D��|�r�2w�!lܜS-f;E'����y@���:�R���q��ϯzt�B	L�i&&��8Y��^�]�T'p��^�z��$t��J�=X[�s; ���H�����F'5��B��Ȳ���S�Uq��P�\N�Q٥�TǗ�[������>y�����~��,�������2�wr��/Ma�9_�[���|P�X8-B:lF��_[�ia)'�IVZ��v�nms���� �7��/���2�y@�VTTdV�����s��bU�M��]��c!nݔ �E��5I�^z�R�K�.b��TC"��R+ɺL_]�h�z�+m�w���3���������9 ��9�o�d��+��� �쐏�����D-����G�N�k�V�P��~� K�p��`��l^0ٞ���%i��l�Q���Q�Yyi���mMf��{yAA���w�R�4i��bg�����n��)��q�����-е}'�I�aJ���昹k]��\4B��-�x��ew��?o�w"B쮉	'H�'@m�y�&m�l����~\!�V�������=Y(;w7&��D`Y�T4֎�Dc����!}[Wr���,�>O����ɣs�S���(���ۦȦ>#��:Ew�~�y��g��jڼl"27r\�󗏿*�6.��p?�"��(�,�[�6�d=���P������h4pN��!�y�����-��,�L��`�6�_�֋f��r
��Y�*q��/���(wW4�����&�B�Ȳ0k��шL�ٿfK7�*oߦ���u���B������@�L�_�޽~:�z^l����P��59� ]F,<�C0Rzi��`,&���x"r(���L�A	�	T�5 A��f�#�M�+ܬX�v��x��y)�����X��y�yX6MJ�ib��6L�<���d��ރ�0	Z���b!;���6���ϻ5F^͟�A�GEG��U�n�	r����oR6�ƪ��LD�`>(���b��w���II�m�����鯘Ab@���s]x`�rb�^ʂ�|V~u�� L��z���V����x�Y�����V|\��NP�+sm��]00��J�E�R,AP�(�]�=4@b��&t֒Pj���8^�ؐ"K6n5��_%;��+�LA,������Ä�8A�6iF���R�K����5P�1@��3�o��݌ƙ�B)�ϐ��>Qo@�d�����{CY�+G=�[�GLAAa��حE��Rc��T}
]�VQ6 ���ߚ;�s-���y5;��{�/��E���Q��h�� $�p�f3�jk�����E����k� 9`p��:��$l@4d�is�2���X&>9w����徔1A���ǯ�#�8?�a`^K�2.�i���@ �6�p5�j�bNOM�|�9�7�P��Y��g��8�ݍꍐN/ᘻ�W�_RR��<AE�N8�l�1fn�oj�o)�c#��'���?g<}���dߠ%B�n�[���W��	�Ф�6i�,/�*w����U��/��6CEF�q�3j]\�Ҍ��ܪՕSf��`�нN�� �F�ޫl666�UC2Z��o�˛�<���ߺRµ��� tg��5��<'�I��Qq�#�`P*m����M[�X �� r�V� )�O������l�KuMM����+3=!@B�Q�S.�q�|��'R"(g�Q��i*��;��;l�K8��������g?EtТ|s-:a���K�*��xU��V�0�0���gǬ"`�и����a���ճ�E������)�,S��Iڭնxg*���?4���� �f���Sw��6�~V#Q����VM��,�vq�|t8����<%`a�X��G(�鬓��2�Ɋx��v}ح4�yt�XvO6S%�ӒJJ���[v�X����S1pC�@�K�9����୏VD#
���߾�������C�7Xl:x����9����1��/��28�u�Ctnۂ��P'[`k6�{S�hw!�h����l��YE�C��HލB�˅�3�TH�g^��cC���7���~�8�n��îJ�8�i�ޝ�$�Ey�R��,�@��y����&�����
:쪒�����qR"�^y�M&YN8����4�q͏C��]n![94�d���q5>����V����^�<B��2 ~���*��zWW�J��ZN�����p�� �����KKK�;��Vl׹a���s�YYYP�@&^�o��Ѻ�]����ޫ��=����4QWW!y�Z9��A��uS �#�R 1��o�����9����CIR�{`��f�4�l�6��R'��l�^v�Q�^E8�k���X�1Ԧ��=<,hx�ʽc���A�����P�jk�1��ڃ�A�<������{�1��*,���gs�������ttt�z�ѥ΢�9�������ſQf�[�n�黻>*@����@�����=9>�.�~��W���i7xh�흝L�*�4 �/6�Һ�0���ϗ/2�%fmEF�:��z�\��ϼ��}/n꧳�������T6�����;N 1����??h�6�.�2O-�Qy�ʃC�*F>O�|����º��K-�g�R��	9Gv|(R�2�!F�#�:��2{ՓrS��aS���I(p dr������Z�󎊊����d�kn�����72y�t!�$���1w�B���w�IF�l4�j/zӹ�����)u+h	��z�X����� �`m��/�+���g�.�R%�]�H�������ۺ���ve�i��jӏ���loKὸ���"z�L�"���A������|�H��.��1�}��Y �yݙ,2݁���4̂tvK���� A"4���%y%��v�}|4ʗb&���Qh�o7�����~ỤJ
K��A"7��#D�_ju��h*�>kʤ��[� ���ci����ԤRM/���ա��Lȕ������s 9�a� ��6���f�Loۼ�*?�Dg	�c*�I���I�_3�6�Ղ�������s��m��h6=w���u ���܇V�a���X͝x>���B����@���ܢ�����B�5�2􈑜�:�y�?�43y�/�\��<����!	d��ϫ�Nc?PXĊR���)� �O������T�׳��ӌ���+���\RbƄk�"�"(˟��K��E����eQ��I�
i�?tq�C)B�;���uo����d�O�2���LSts��ؙ*Q�E��W�?��Tf;�W: ��q��Xl}=+={$˃*;Fȝ�*S"��x��.������XkH�픗�w&�J ��x���g���f)��a$�wG��>��A��^�}�|��"#��z>�LW%���$.H���S�cFӤ����]�1�on�p�9*ZJ��6�/7:��}��HO��Q�^o����R�l�[���v)��g��6d�0vO��F�[}y�;�F��C��A�s"�l����K�v�f���{v���h���K���v�C����\�}��F�bI���f%�:�{{�
�L%Ʊ>�{�C�}|R޽{�.�E�ͬ�=�Ī��Ē��e���u-��1��nX�Q��]�h�}�؛Y��|[v!����Q�ˊ���g��:�#jN.Z����ᣒi������^�����9(ం���\��4:'�0���,�~�{��@�m'GV����׹s���?d*���q)>�2
!	�e���ܳ���A��;��Ж[���!K���᥈B=���ez~�z2~.%�y���X�������	=	~g���k'�r(y��VLH����ݠg�����d�O <�Y~J�n��W(��h���v��=�ⶎ�+�p"C`+�G�vy�k

�dn>>�Ý?~�}��5M�[�|��ș���Xrh��$�-��6H�0�4��s||��]Ĝ�_6�|?�D��5G�DV�%��&}�S�D����ZtDY�*�ߤ�x��g�T��SXk�DL�6���9p���v6�������4�$��,�-�]���E,C�(��c�J��u9Taߓ�'H*o[$��P�f�`f�{�@�B�T��NT�j��:oN7Bk0�N�	=����S�ר��[�� �X.�.�:��r�f)K����G���p����ǖ�s���|�k-�ئ���P�_�ʀ	�
?�T�}��%���Gm#��^W4�j�e� u��=��5h��h.5].�条�df��������!@���RC�$�Chjv�
�o�>��P�n��s+��3D������²��Q��!y�2��sՙ�H�TYp��LΌ�g+e���;�+#�i䨕8=I~pBz�1���Y�}��tû���G��$��z���I{zv�:��&zE��h��$���-Ռ���x5��	����
���QQЉ&ҝ�x���W=0���nԝ�ݪ����,��Ʋ<��i�#��B�����[|^ԃ�����<ЈGi:P� ��q���{�$oܨ"��l��9������(^�nrO3�hyKRA��tc��W�w*�R"��@B�EY6�Ю�N��,n��H������A�/���(�r	if�r�P�X����Zw��6�p`�j�*#	a�S�3��N�ц��X/	��?d�CʒC�no�/G-/�"��"���Z�z�$q��+��~=yv+Q�&�=�9 -��s�C����wC��0��c?�Y1��Ձh�����i�c>^Պ\#�Ta3����"3��v|oCd,+�@D�����Tn^����n����Cw�CS���Uk?Gߴ������EN�@Z�ﹲ�(�z��:u:�� �NA�js�q�F�@ΐ����Y�E����8��0����y�UiJ&III}¢���իW�!䝯�}���m�#?�$�oA��	�F��z�̴���z��(����������&���N�s����M�5j^Ck�>��]�M��;���E�~}~��m�Yh?�#�7�%�;qU����g�է!h<d���N7��u��p��,�*mCł���	E�]���'j��{7胸0p�j��8�iEI��w�E�K��Y�7v	f%)��֟a�7o� �g��"�|��Y��7^�<./_h�%����L#p�_�Y�g0�lfG��l׌+�G�{�	"��u����q�-Є6�sr|�ZX�Ub[8*{,�~Be�� 
*֞�+x�N<�xL��Jx�@�����?ڭ�qZp{�D�籋�C���/\�����NY�掣�K��x���zү�X��Ú�u���%)y��[>?j,Y+|NԮ1c�.;��������j���y �9&|~���:wkѯ_�����z�0;�Uyu��4C����٥h&�9`��xAe4�m��/?�Z�C�����tm�]�J��i�mt��{�3� �o��h9׶�Z�9��H֪��l��s��#��"Q��B3w��2Y�xH����0J�K1�����׼�ѫ�F� e��1e�����W�����.RO���G���؞SRQ�k#M ���|�s|�s��p���jzSJ���0��T�����2��ow��H���?�(�1�.p>����KX�J�!�r��D��ۑ�r�?-�l�0K1�o�*t�[��|����&_����Fq�/.��k��g�U��Z�M�������H�r������A�m�=��� �x��$+�]�
�v���XQ$�
�xLSN2Of�b�|)g�����{���ljt�������d�YI�#[%`]�:��S�F��~��p��y=9��#�n��Wh~2��
$ag����hĭv&@^�"��g����b�&bd�͖q;2����0Y���%=H�v����|�G
�a��|W+���r�>�)3.s���{��_���>f����Ĺ�K����˨L5n�*X!�Sr���y���\�7����!���ͨ5�5��}��z|<ʍ��Â��E/٠��V�%����8��"�$$��{���x;8|�8�ݕ���-Z��c?�����V���K����e��\�����bh�X�b':n��{���@�C���=O�|�G[b�0�LM[�͉�u�"��缊>\��9�q��s�1��ZI������֤4\"
G��g����,�����&1-Qu��@���;�'MTy�g㗻��:�����/�k��qo� �p~�,��N�ҕ0�G�s��q����ˣa ����
�c���}���٦6��p��Ԫ춪�]k4b�"������sR+�0��c7�������}rX:��p�.ۓ�T�w����+����ml�3�CyRW��wZ{d�E���z�����RUUU7����N������j�5��ku��u����	���)|eR;�6��f�s�˅eS6���f�����
D��+`�+2�l6��-4�J˟
��fc���H�¿�i&��߳!�db���+�=Ey#����Ua`clO>O�.�)��M4+�X�*����`v�����E*�.;�����;�ئ^(���l��������5�pE����)I��pU�;n������lpne��%*�sxW�u|`�D��xh}0J��Q?~�y4"�a�m��<��e=��j31��?j��U���_�6�0C �o���~:������-�>Xai�h?� ���*�j���b:/ܻ����~]~AA���������08��Ԛ�w�ט7�1�|��ND���	���o��s��m9?h�ݔ]8��d��F�Q��4l��ND��~V�~���x+�8�>/����
�Y]	��V�֍x���Ǚ�~��,g䊗��8sN�r��F�����$:Cs��n���N�G��S�����r羱	��H�WWW�=�	����)�f�k	���Lr^Ц%U_1�F'���s[q5��P���|�O�һ[�xP�a�C��Bȵ0_#��Ȍ$^qm��S����o?�p2 ۮ^�[};�կa2m<��y�hi:�x%[��2RX+�}�`�`������e�a��/#V�be�Gk�^�	</�]����Y9�ؾ��{��;���DWc��B��E�C?��R�L	&�h��H��t='���РsE�PHP���4�`��8f����7��������[g�};��.����Lك��C�4�E�x��Q']D��^���lN7f)b@6s�Z�@��܎�/.kJi$x[�/&GR�@$����߭�#<�%ݭi�t�E�R��@��@�dĊґ�;/Q�S�����!L~�c�l�8N�z9� :"�R�-�W���I�ȷ�("��[��BBq6�A�@G���j~����~Z���-E�]��79�o��_��c
�t,
��fV�8�>�4���9��o"?�:Z5�l�������{\��?�"c��Z�I��6�ZS���R�ڃ��5�!-��O��;��T�Q�f��P��M���ڳ�拶��^P7�$H#����z�_�X�6�!c�ea"�H��A�w2QW��G )G3l݇(	�Z�X	��|��V��=��d��q��XP���gk���r�΄(�Z��?b4*�_��$�֮��U����I��-�8�#���:��N��u�=��}\4F ׬�Ѽ� ���П|���g$������/�:Uc��%���-���e�v���5Z�lJk�X'8r����^��Z;!�����N����l���42���1AQ-4�ט�\���O����d�h,����+��D��\'�#�����n���(�Rcx0l~b�1�6:׻x�0�Z&p�t�>-I����{���:^�Ȱ��JD9��5]�D�Xo���ײ��Ƽ�:b5����I��{�ܦy	��T�����������V<ؼ��$���3��rW;��ɔ��̥���R���5w�4�hDz�gGCI|�m'��[[{�b�+��22�q��?����n�O>>�Q��3��G�;5$�z�ދ:��WyZ��8�lA{�M���ɏy�w�����-]/� 'h�/�[�o^����4F$ �^Gn��`�u#�ZkS���_��Ϩ=�Qjڞ��mGVh�f�]6?�kI�N5����l�E�M�����=ڏD~%G�H��3*�ݺӤ�"�I`��'k�����GݾM[kC$�]����??�#�����ǚ%�rR}��)2���i��۫'0�r���q�ޟv���#{<������C��FC�돣�d�;��|��7P���oV�X�f�A��#Y�ץ�rD�-L�?y�PT���7F����7���R��/�x*R՜[��O�0��g9HY������*������"�9)����T����כ���BI��ͨǄ���F�'vɿ���04�m���:h#F�d��"�O)$`b�MI1��*�/L�0l]�������w=����]��*R�A����e;����Va*�@�`n�!\��%S�l o���0~�'�\ �v�n���	M6��t�U1}�қ�7OR3�S�4�v3��?a�c�y;{~�B��j{�Wn��ã��s�{H�u���PAm�_���ٽ����8�Yrd�ng��ApwJ~���fsZidܲy�)��\�E�a��dl0�4R�tE,�4ƚ�0�x�E>�>��wK*)5�-���K1w}���EҚV�k���LK~rzo��,f�[��9�Vd�ћ�☆\��G;�?$Pj���hT����R�c�z�D��a�u|����M u��=�]����?�0 $U�h��N���~�%�[KU'���L^Q��% ����+�ϯ+`��pho֚��_��fG#L�luv�sc-P�+H�Σ���g��ϫ��	
�#��4aUKWD"O��ޛ<m��3�U��	��Af���2P���Ғ��E�~��Z ����hī�xω����=/3��6X�WO_ެ�� ��Q�8�e/�F�D8�=��c�J��N��TOꆞ''(�D}��R��"��r� ��w儜�F��Z���mRC��/��t�2��T@�`��˻e�9��@N^��K�.z:�V�Fj>�6w>5x8�S�k�Ba�t��G�2FD#��Za�>�L����s-qF�sa�?H�%K�wM�6�Y������	���.-t��>=�iR�C,f��wc���wt�UO��9M�t)LR̓m3����+l/S	�<6�s��)>������{�\���Aq�_�7EAS;ܱ���WL$ztC�?���ID�+��!�+�bHV��N!�LdIp��Ǭ1j T���#ԯ���6����_.g4[��4}#i�v�ߞ=�&%+t�Aώ�I	�2N����'�[����R+���;���h�X��;�[^5���Z	�M�mMM��P�Z������� ��9 ����������Q%���|}�ǀ�c?i����lNg:�ɳ*�~��0bc��lVE�l��l �B�[�'H+_5�'�.��B�����[7�kEH����K�}�t����؝��Ȥ Qc`~�7�E?��IYy�� �ֻ�5ZaCK�t��i�`�gv�N}kkk]Ss�N���{�Zu��N�*+^5f�Msh�g�|8����M�2��_=e!�;���ɸlv�7��_��v��M�(|�6k�X�2����n/*� #���eT:k�"�wp�p�'VM�6����0�J���۵�]%2/�&�^�:E6��E��T�#�]F�{�1fi�@:����>�vU9������jqϲZ�/���<������h�qq����n��%rM�j�۪ ������88-S���C�D��j���T@��sJ�7�O���,0҇��!����zP���rр�٤{��l�ھ�T;�T�!:��/�<J��&��i��-T�r*?~�W;RoN�Z۞^`�4fd�[�N#����1H��/�g�qթ�9Ȥ� �L�&ZP�\������#����5�:�o.�&��4�$�ioQT�X��B�¤��~=\2cgO.�*^�X��I!����S������+��ܹ�y� �ޟ/4b�n(�$š�?рiL#�ؤ���RG� pQ�8���ı/"��KG76���"l �	z�g��Эq�UV��?dX3�%��
>�>�,_c�)�}�
t����D�4)2��7zN��X���?�N&��s.!�����'���
bx'oH��6,��N��G8�(�&)��q�)~4r���qO:j�PB�i�&�L_���?���. ��d5+���t�Z���o�Qٵ�����/;��ݴoo�GG7,I��L@K�S)�֫���r�>�����������V7�\�[1R�c�z�A<mS�k��~��א8��,�,P-�7p�T|Ƕ5W]k)������PΣ�ū���\)��`��Q��=(�cNZR���p����p��! ���~L2��/��M�������Z����QjUgV�@��ٟ��"q�U�U�^�ۮ�m����B�f���|��=�-����	�M}	�.x1�{O9��L����y>ZB�R��Ô��F'�B{�
Z�v�NP�s�t������_���.ȩ�� P��#>���_�]����>��ʿ�q����/Oy@��x�4��="��_	BK5p��v#��,���h��4������=�F��S�Aۿ�p�*,�������'��p��#�H%AowS>�r5B��L������z�W����gg�e 
��s{���r��Kk�����HV՞K:>�Iz\�������wYY�c.��G�������]��)&���T�9N8!��/R?�H��17tK�+�1�5�.�Oc�E�Yr-�',��Ts�����C`���nl��C�~]Sk&p��c?�Z:Dp���U!��ۇ�8H9��x�c����%i7F��d�<�ڹ�Y|�0迎D7hu���,},�@�_����%�!l(A,zz�(Tm�b ��5@��Y2�bx��4�"fMi����)�,B������`�|��ޞ���(��� z�8m�F�{̭��vOi;z�����Z�.:�z!��R#����o�������JO�s-�n0�Թ�C��}�y��9!�g8�+������dwVmuꯜ�q��jsq�qs����X2�{8@�5z��Ub8.J�!1W�B��"z=-R"+}�]Г�V���q��A QVv��ڪM�@
VH6��,*�KO�8䴳(�^
��XU�r`}4��ϫK�__��Ъ�ӿJ�:���^�p���:�
�?g.
�}��þ�~�)�_�	�V�QٰcG V�*� ���T�2�F$,�>H�h�Ӏ`v W�]��l�]�
��m@r��m��hzJm��#\�����S<g��/z��[��H������ɺ�LE_J����|�g��ƌ�A7�ھ��V�g�Nו��� �ˬ�t�WЦm�3l&�)]�h���t�3�D+}���%�gM�f�]q���j?�~�ދȣ�cX��8��w�n�PfPt�|��%�sy�:�N	����"ܻ�L�S�#pԜ��އ5�,�O�O� FH����T�[��
����	P��I����$��T���x@嚕����ӧ���z�'�Z�&��~�z0a��t@�9[�%G��Q���r���b!��D�-[Q`���'4~ld�S}_��L`��<�����[��a�W�Ŧ��Οģ/ځNh��Z�p(X|1��8s�Zx �-�A�x�ʝ1o�t�ʿ[��\C�ҩ�\� r�K�hPuu�������eĩFDB��R	N����,� �\�}O@���������"�F����O��.E3��pG��)��s��Ȅ��P��Or�\�3ۀ�g	d�[�Ag���U�hE�����R|I>�~ŵ	�߸��ٲ��7n�5���fd��X���O���D{���5\�G �klBp��Mv ���r��? ��C��(�J����)d����BP)�U�y�C 7F(�����g(ݨBN��=�ѹK{�5�7S�g6�_7��~�rp�J�f� ATj��
%7,IK����Veh�r�a��<�p����d{�d{���/�M��c��m�~ ; tE�tp�돣N[�p�u���a,ep��	��t~Z|������I1�s��������\d,�N�HZ��W6묆d&r�HhѤX�|T�/��vPk'lS�?���	l�K�"�X$P�c�%RtM�&��c�W�8�ٔA��$Z�Y%����4��	[^�]L����Ԇ��џ�vw_sQ�����y'{���^�.fp�Ŕ�"6�}�liX���j���v�+����8H]͂Y��>����ĢTiJ��	���g)6)}�B+�߿ �04-^ı,BO#I�PPP��ugUh����r�t�y�/-���h���l�ٸ������3�3ᵅ�a�d۷��h�;:�2Z}��aq<sXq��귌�?��Je�`���M�vI�B%�M./;L�mM��7`3������5~������f�͚0�g="��4ʧ\Dr[��Y�[��O�ݹ�˴�P;����_��>��RO�ٔ�bX�� �*�=��p��p|��'�k�'P���̾{ �6����ݻw�0��U�[;��{�㘋~وA܆����m���ǽl.cT�c�@��.ES��9wk��g�2K�d���J��Q�z��!,jR�_GA��;��;UJ
 
��ƈR.]��?�g��/S���A��C�#Nd�Olx v���a�h$�����_�H«(*���Ř�K���D�-L��{�b�[>D�ӝN��a=��F"���^&$���C,0�կ�����[���/��V5��T_o�����FĿ�8�� &�@��bPw[�������i��eh�A�4�N���T������}[�tS��Ѩ��x�Ъ�e!�<rؒ����E��'3����ǧ<�%�/>�p��]iz��7M�1~v{r΢���И��Ŕ\�����lU�����B#9fn���s+������tz?(���p��`�3�n^�]�Oүç��=L��?�خ!(`�=\j�I����A��)�ޚA !�X�eZȾt��1aͰb�S�ܠ�3�zI(�ԓ�仢���:5h���J�$�(H9G����HX�g�434�A�,lk�*�5|?�"��<ʬQP�y{���$��45���3Yvf X2����Z]B>��~l}��p�	J��-Κ�'P@
B$�rn�y���Y��~[;�����~���y�̃׬��rJ"gb��D�9+����KY�_(��V��ڔ�.R].�.�Z!8���ݘ��`C�S�z)���>��ٽ�%?��jn8AD���״���-]�ZX���~. *m�NS*��,za�O.��&h���W ̣������R˚�L�u��oA�Nc�� �K�M�/�O����64yL���n�.[�D2ڬ�͈���S�j� ��y<w���)��}�.������=҄$D�Rd�ԉ"߼L6����c���|!��\�費A�4�rڎ-�Ct,�ct�y �k���R!cT�|��蟶��E���XR$��@R
�#έw�.���E\#���4gbv*.z�Rc�T7홏��I�د#nt�����?h�=�,b3NN�l����c	6�׼M>������Q�	.���SK��x	�a<B�E.�Z�]s�Z���߈��� 1��֐�D�=S������T����V2Zf����H[���ZE��\�"ԕ�F\{��}�E�-���е�_o�����N������|�����B�T�����Z��KS���<�?�3���%K�V�A���+z�Ϥ�q.Q��':��?�ُ�=�׿��84>ZA�.&�
��Lw�!\=�3�=��'Xc�$AЙ�%����1�ָ����^���7.w�d���C�),��I.qʐ����{߯�c ��p��ҝ dj|�a�� ��B����Ʒ#��~��}gy�oqg7�C�ڌa�m͡�ÁB^y����dv�;��i4�5��]�\~!��Q����<p]žEc��>���P���c৞���4�8��̸�-����L2����f�;t+󉦔��F��l�dK����,�ݡ�c�pg�E�iR���#T�/��ۑ���fQ�)�߈g�����^6�3����!�bE~�&��ş��X�ؼOkג?�����73>�����
Z���u��{�旆!�������oP�ܦ�j��0���|)l��S'`S�P��?�S_s�p��J���9����d[�T��,�Y�Е�{�QW����<�G\��,4�i8l�A��͢��Tm4�C��3�P�$���g�CE28}��З}�tZ,�L_%�~�Qټ��]�F�cv"T_�:
5�օ٬0j��S��m( ���1���61���2�)�৮@>|�	X�[51��;XSwy�QG��\a�u�?ſà���Gg��& �f�Z�% �Sg	�`B������9Ȇ�Ш�X���7��x�d�	�n���!��o&�P.��.�ڮ���e��
��K���G�	�~V��}2*c�UC|Z��Y�����B��$��F�5 ����7x�jEct��݀�l�U$]��{���"]5�~���B]#4��acN:V��OZ֊L���ts�Fi����5���	z8�N���4��2RLD����1�u��~�����{��f���,;w������Y.��aX���bE��������F+��n]�/5�����>y�[G�z�J��f�!6/|5iv���h��Ȇhሃ�;4�#�}�������������Fb��%;��DI9��,��ڧ��v��]�,�z�)s�97 2����DLQ�dKl�U��9!HoI��ܓ��J�.����E��ܜ�[���T��{�E9�c�����W��k&�/�CշEA���=�%W����_.I�s%��~�7 \�:x\�|d�U���W����c�ey����'K�._����B���/b�����E�^O�F���"ԗ�"�� ������>��h��
]. ��ؕX�H�9�E~)z�ցb��0��&�LŹ����_2����\y*������W��������JQ��dpvr��S$�,I!���r��띾�h�&`D���&�;�i�J3����F2jcû;��Žėc	�>g�c�ZZ9��O�Ζ���5Ł(���T�|����`B�`*9�D��7
h�������1�/I�e��4(�$b2�6�k�]���:�y��@wN���B�f�ϒ�>�(a���>W�=��x����R�A�{8�3�����/�C~�4:
�8�^ӈ���}��:c3����>�"�-��ZhKЉ8+r=fj3b C3}�_����b��c�ae�Q'w�2�BefJGcP�c�m��Pz�q.t��`�%׼c_;��?�]���q���{"�wHE3�VO~(�|3�~�j����.���g�x�*��*,G7���3��q	/�Z�:� �uh9fA�Yb����@*S>F���>:<�i�X�I�-���W�����/��>׸Ys�S��7�7Ug@����h�SrJ���袅����!���>�&��M(�7>����l�^�H3z��sj��g������;��,4_p�DW'g��;Vfl�t��|_[.%�m?/d�?���8J7Tor=8@:�2(~�(�R�W� u(	���W	�Ǯ����`n\<p��B�
�-��~[㪙��s�`���]o��$7��O�v�G�<;h0��^���S�_)1���>�u����&�+��e,�R4�:�Eȓ��W
��O��$���̠,D$x|3~�~+�/ ���ac��$R.�:�
p�7�ǲn*�:�����i4Zjb��k��rJ�:�>o��R�U��hdl"�P� h= 5�k_�f��A�6TJ��	��R:4�s��ZvO���M����K��5��O��3`�X�y�y��	��I9"^�E�Կ��x�g��@,(L:��,*�n��s�$���O��$ʓ/��
���2O���=S=�BmBr�a�!Q�?�n	�٨h���������<(�x�~G��0)a���bXu1��p���"g���R '��������E#����=���**aE��O�����~6ό���׀�u&�=�и�<`�գ1����_;�)Bc�}���Э�~W�)I�O�a�,5*�*,1�1��a���_��'�I!N�Ms�f���ޙO�;v�-�p�?SL � t���U��H����\�e'O��%�H�E7��#E��H#�+�>��ܿ�cH�j4��cȴ1(�
�°�t�)z��;P@5=�H�?0y�$b>�)&�S 29��`t��`K�T�bqhss�}���F����|{N��p��r��L����L��f�:;��sB���u�����,�E����+���z,5Z�m�Q7��\��}�e�B&�0'���p��-N&�(�l����?&��āl<Q���5��c����i��w*��iSrf�wMxI��UN���W>�s��� .�"
O�d8w��er+����rJ�R)�����1¶I>�D�8�<X���:�_5IIո@����1sS|I;6�RDq�: )�,�3m�p9'x14�#���ƑOY'��!�9t�5z��5"F�!�����;����c�9M�wt�����8F��;Y6~����J9� �BY7t�+����lY�m^8�p�,��E��X�d����x�u[4�7�8�
h���"���� �{��w,,�;���r#�S61$*c��IP�

��И��q%��Q�$���`__��X��a
�M�ad&$��ᑃUd4�c��9��A���{I�;�����ѐ��$+��@������v�.����&?đ0�@�e= kj_m�����xX"t��$���bݑ^�"��������@�+%�Z�/�?mѨ�֝�&;u⡦�͔�{�=9CE ��
�Ñ�K�@�@ɻn��X��R�t4��L�zG`�ba��D�S��w!���^vݤcoBW�(3tX������Rʬ���Î�^���JGޞ<Q��s��e�9��$1I���PRTU�{d�����7�[�˷�y?Փ�|�I�XF�޹j\m!H1x_8R����&��N4��U�"`�>%�Et4X&��G����{�w[���}z�
k{]�[�{�0^/��u�[-L~B�:1�;m�\�IkO��^��@s�"�p=�*@u��'��M�˙F���C��d\�]L7	qp�}|�{��1/��'�G�CtF�ߪ�L-w�}���l��%���^J^�ey��z,N\\��|N�i�WT��Β;����B�T�e���k
���!"�P	r��vbV�yu�_�]h�%��K�m�f�����Lx\xZZR}m63`|�J-9�r�N����l�{^�9:��U����i©�'�<�c��"i�<�,`�oѦ��ﲗ�y���Nw�Hɾ�9:��}ΊH��p�H6&��54ۦ�_9"����+����t�l�x�ĭ9pp�J{�}�p^�{���J_2������/P÷�
������ ���5�!s�:!��l��'�L6s8�*=bʬh(��ur)��$O/�H[z���C�>X+�Q��gX?�E�z�^櫳���`:�38�(�r ���T4����?�P4���3a�!�K�e_��m��2ƅ\Q`{����wq#�o�������T���w���WS��(�h�QqoT�@K(1J ��&Fp���`8I[�I;i�8
L�K��~ʀj��ݻ�\WJ|�V�/����}����K� �"oh�SH����_%�Ţ�B�v����w��7��c��6�ׯ�c�F��۝"01�b���"���B���Ξ������.txoj\3��ãz�O�hB���qYG���{��(��d__�$�����ih�F�l60���U�8׸�F�!/N�PM�����G����@�o�2�<	=ᾙt�6|�8G��z8�v5&���(�ިq�⥠���N߹�&�&J����:;!����Q[7�)���(��y��

&������A��]�3@W�Og0����
���J�-$v�B3~b�2b�|��i�N����,j��ǩ�����w��0����&��L^$;��
ੑr��D���dQ�S�+ާzUu��S^�?��]�@?�Ky��*���4H�L�8�	f8[jp�B�/~������.>���b����|"���q�.�5{������^�'��	���m`��jz=���-�x�*z���۟gd?q,��#�X��(|$�p0U?��-�g���E{����er1h�?%*�H�?B�-�GS����]Q�/_�GU܆nA*����;W���Ls���!$���C9ڱ_������"O�U�H�& �?�=�_
���\�zd�A�)��㗝	��7Oz�:��׍��3�vjJ�w�z���ئ?F��kl504�e��{�W�sK%AӉ�F�ŝ��w���ûζ.�����D6[�!C)�^�1"S���L�#�`���hm�荛�Z
1bv38��B��>n�}�(q�TQaoc�+t'<��ߣy������/����:텒�Tg)h޽�p�� w�=�K��7ۗk8e�@J�"�$,�&���=�u�{�tc�7fzG?���ֱ��j٠�w���j{�Y�kO����%8*w����<GR�n��hc�n���T�/�W�^U�A�h·3�*T �TK����W?��J5���D��� _�E�{�'8v����	��&���dI9:'��As���^���(�Sm��]q	H�#�]����!�
��_���ip�B���ÝUA�v��,��~$��aa������9����_8����/ۧ�������_?�o:�|���ၽ��2?8�C����	�}x�i:[��y���0;�$��'���GSߥ�Ε�����/�w����<C)�g�*Vy�����c�gy��ˢ��dgUSc9� dB�2�۫��R�ˀ?��(E����m�V�st�uZڝ�P4������_X�N��(z�MY�sM� ]�,����$���$�����:{;�UC؞�s��e�Q)$��.�8K�7
��=47Ϡ�憊t��|��E�=?�����KZ*�=	�ޠ�s�:��l1���R����bj��T�>��C����ZJ!����]o���(��"�_�|B�ك�����G!�+f@T9�l����A��� C"��N@���9x� ����l,�����J�0��������$������w������H�{l�,�e%�L꽯8LR__ߨʈ�̚\a`9�Z���c<DBkk~����=Ѓ��s�%�=��=��M�U$�W��/�^���-��2�v��u�)�)��?�Ru^"�Ǭ'��#[�:;M]�Z��kh��������7������Z9��ٗ�De����N�'x�*��^�~a�����f~|V�+��řw]������Sg�ST�vZͬA�&әq�*�%��T�vxx�a�֏~���D���v�S�`�ꂆ=��6���_?�����W����H�h�Ba�����!���4{"ۊ�i�4~J��+en2��Ěf͋>�S3�� �j����iF�	�hP�H��-j�oZ2���1\#���N�M��l�]X���$̘���u��7����&o��]��n�^f\(~q��֘?�����ؚ��������)�UiQJ2Qq{O�0'C_�X�NO8j��1����A!
O0��A[Z�\Z͔`V�>Kj�/��(�E��bȖ����MD�S���K�Ey���b���VE~v1q���歳`�*w�oZ��Y��߼m�Pv�P"_�x�n/j�=N+�5����ϟ༸q�Gc��pt�z^�lR�,:99i����tdk'l?AA���Q{��wТ� �F�.��>t��^Ԅ0#��h�I�`���r��7F2���G����[MM\����#Y�d���|p�4t:�5P[8%�'�P&U�vC[�B�N�)&o|��&&&B�@��GB�<��Y��;�iM'$��,bo���MXCa�t�!X���0
WuA��s|L�G��Ci���^8v���Q����4���5�i�`/2���	<��SE;t�C��D�@����4�U=l��z��Аe!)Ŕ�"C���P��@��s~]M8Z��qw���o$���0a��go�׏#�s~��N$��"N�b�uH�x��CӦ�/�F�j�У-EEE���<�U��ΉY�R��;��c�����
߉���_OXoŻ��(~j��5#x���;CΜ��;¢P�9ă�2����_P��X]]���}�뇡V�o���D܍ T��|�����ih��0-��
�6ι@7��5�!Q�#5�~x���w�l��y�꟏����ە����(__��������j�%q�y,4��nTO(Yh��o���/�㷭���f��{�>ڛ*}��l^↝�h1�|���O�K_��]#))R�Ss�����}7O��,�j�/[/6p�P1;w�s�1⛶Q;��lS6޵0�?�}o`p�>�F�����N��88^>�-�[Oh��+)�k,��MD�ׇ�I�S
`�,�T��nJ��+��|yMM��DJ��j����� J������ǀ��� �O7Wr��!�8�69C�?ws��~�����&�Uό����3�/�Mĕ �i2�m�p�z��2�3�A�J�F
+�B��D)�ǿgS�e!���$�L���Ϧ�{���R�d�7p�Q��LM1M�]�:���k��#����[�܉��V��K/(�ry��`V�F�l����ki�Έ� և�D�zf��!��GM���}�!��'/��K�<�˚�A=�q�i��ё�H�:���h�14�7?m�,2/�_Z"W8���X4Λ��Ѥ�ݺ,�;�u���$��=U�L���N����7�I���V���o��af�,*H��m��q�\��ntM)c��#˕�L���w�gk�J9"�p���g�m���$Hީ�y6�  e��W^_��ӆ���*R/o�7���LS�J队���T��_�A���*�|�>e��yۗ�cT�X�
�f�o]�N��N>V֮��˗G��Iզр������(u�2*i�w�|
�R��s���P2
�f���̑Y�8��KY֛�
;}ӫ���_u%r�H#v7�-|��1���V�1��T���3�&S����-��~����[4o�zz�n�rwwO�����ո0�Omqx����~�Z;��:�Ȃϻ�ƅ�;�����I���[���5�1�R{<�9���~¬�0,<q�{� ���jd��W"F��t�2�z���^���7�*AF�k��zt赙	5I�� 
�M��'-,|h���,B�\iԱ��nuR#�͂Ỵ�-�#��8
Mu�'?�:kk?Yr���P>;�I��U��� ���a��Io>G�ڙW�5��՜�6� �N�k�h,��W�m������	xإ�2���7%��D�+a�"Qd/�;�x�3��O�c�7�O�GAՐWP��"���ق_�/�^�)�g^��!�OL4ϯ�Ȟ8��%ti�"�t�c�f��&mn�Es{�b� bK<S=� IG��jהOm֗�KZS�20���<{�:�h��(R�~��1�N.f<u=��b���)�W���_mFpݩk{��B���ua�~Gm?��n��K�t��A�I�������림j��&8�"8R�;�[�n_�L*ICS�%��~?<|������0���6���R:���qN�Hd��`�� �}�y�Gt7������D,5Y�8(�2�_[�B�W3�8���}8��|��#h�Y g����`d:KA���p��N˦��0�ε�~�6��jm1ֲ)�[k.�%Ś!�fJ��3c���tC�FFF��m� ���B�N��Rf?rd��TG����)�����M�D�H�.�s����A�qXx�Z"��ن��Q�w�ɐ~4�`�G�n�ӑ��1�~�<��Z9�|��37B���b@(;�Y��x��;������mL&��k]U��\�媦�F��s�20�����g-N�x����6�;�p��`���D���D�n������L�h6[7�Ά3�l��q>8�g�c*��J��ۚw�$>)���?������}�"�h�O��0�ą�
��N�cy�L�ΕH�� ���?@+K�|c�|�2<A���Z�G�тn�ZKu|�ds��E$�U�a��8]C+�2���p�����5���������E�sqX���7��!5��g%�{>|�.���#<��A��*-vzEO%~n|��w��i%��&���T�:�'_�A#5
Ŷ�{�����m�[.���������{�y A;�׃4�V��`�0�C�m-u��z1&rf*v�|k4?�zGcp��]����@�4��zg�\�������6�{DN�v,I�^Ki�aV�G�Ld������S^�� 5Qvt�o���+4%}=f�K�g�������7�൪p{v�%�瞱Ǭq�8�&���\o�UR����~���QƗe�[f�����RQJۺ	��S�a�JŏVIۯo4�$�)[vg����6?�Z�s�y�޿}L�!k:����o,]Vg�����<���q��ӬϰDlm~�m�J�Xm)��Q"���+w��9x�Q2��xskk/�壍huv�t0X��R�[
�>����-�a7�Q��ϴ#�h�� �k|�M�WSS�WǽX���'%���_&�.^��+���kk���>���g�d�~�鹸�FKٔ{�8�[�L��l{���47����5�yB���V�ꟗ���D�;�$t���/n7�+����9xvѩl��(�����2+��%L�џ�J�K�A�*�ڤ�_��6���=����[O�b�&��ws�m���"��M�� ��#��n	�d�:2~fN]�фh	��P���p!����j\B)���!��B���9]������O�ɚ-o����_go�Ā�	H�J�P�>I�/�q4�Q���!����Ё���ul�FU)jس��q~#�[��]�'���<mV|a��/����eW4z5���(�n٧V��T��ߴ��^�i�/�^�EG]��G���޹N�~�b�K���M�5��n�o ��7�_Mp�E$�6�c!ͅ][�n���JW��^�P�B.@9���e\� �A�6��Z�K�x���b�MsGqx�:���k����ƒ��h��
n_��`���qr�PwL�m��R�Cy
�tJS�"�ym7?r{d�t�ٻ.-@�:�����������,�7B���$��9�u����X�X�Jyn,�ߚ�1|������5#N������5KLϥ�e'�mb�t��^��Sm�۰�[���[���]�����U/�BSc<*߄��T����om�s��\dd��D�����R��=m��#�q�Z�����n+�����e�L�_�Q����dk�b��+�-����H��X�ۙ2�����ȭ�yU%����t��Qz��*��],� ?ou���^���Bn]��1h9��T��D����I׆��wC�Dlv������s��sن/J��0�fz�I�=��Ԫ��G���(TH1��)Zh#kt�R�`�4� qxtѩ���#��2��=�E<���s� `tE�>	���fӞ�y��'�΄\z�&��Z~t�+�ўX�|Q�/��l��D_Vh��X�S�i<;��l���l]��97?P���r:�C�_j@�Ve��ȅ��o��ثu���R�ᯚ6~�6=�җޫT�U��af8�����~_!.n� ѤN�S���w�8�y�m=� �rۮ�YS��:W� ��-��F�$��D�]��7N"n������`��M,�Y6Wۻ�Ԣ���sEI3����oztˆ��ԕ@����g��6��h�>�n\BiZ@}|���
����vvBs��w�#�`B�v� 4-���7%Ƣ`�����{,��V�{��rW��}2<@$o����:Ԁ�����"X���z���\�CYF�+TI:�Դ��O�����G�M�2��u8�v�|j�H��!���?�d��}�O0Fl����=:�G�}�C�){���ѐa�,MJ�Q����2�v��P=����R�����ϗ"}�L������!4��`oME�S�a�[��y*��G긮}.Fh���^桇��&���W�աz:;���K|9���#��1�k����Ҥl�>K���=����j'n���|q�/�bX�ܛ�l�QQ�۷/������tR����1�+��ܪ"��r󡎀��|�����*��٧��	�I�k=�V:��!���]p�kN a��$<�-:��r��#R(e-�gI�
�AIiiO��qO��"�:���x�!߸�ܱmm�'�˔F0�yw+(����~fy������[kZ���n�5�_:��]<<�i���哪L��.�v���\�����[*&Ĕ[���{g�An��Tp?A��W4�g�Ζ0r̋\J\B�����|���7���7����_n���O^�Z��\�L�.J
3��N���aI�;!0in�Va���{��&�����K(�0gd4��|�h:��k�K@�O�d�m��J���h����ʎ�3�l��ZӃ��WV��P5��xئ@ڙ��*v\��gN�g��1 x&�F��'��aE�Vyj�{���>5%�3�vٻ����{`�-N�)d���}꣬m]��P�i�V��<p;�񿴟|������b��usrz�3'�զZ�xH���&�ێ����V����H�����V6�w��x���S��S{j�?�ȼ�_�}Ɣ{��a��yf�M:d)v-:ￛx�Q���*Pp#J��������Q!��V���w��9O�4ϖ���1�>D�S/�����]�������H�%�>]���b��J�[Y�ۥ�sN1�����ݨ�/&0L�sy����/�^�	����*����֪}t�5�]㯉��ޱ��Ah\���ݶf+�3'�bemYEr�� ci�^tdѕ7l0D;o��vi��w��&�T��t!�p5k�K$�د���4ߕ�Ȇ��x�/*���/�����!sDg���~|���ƍ�/f�	a��^j��SiD�J��p+�^�		W��(��Pk��Ly���+[`#{6I���%U�r���R�/o�%vQ��Z/lv1��Q�`�Qv�J�hsrNj�Ϟ2�ц����y�W�c�և2,�K�;F+nʔ{�2J

��3�Hc	�R��$G�BF�n��ϓ	�AO?��.��N\ӶT�y"z?a�м���ߊo�@������~m��a&�b�����[+t�:����@���8�3�����@�#����{8��n�TJ��XbxR���?!�+nIl��1�����wG5�@��uTT��4P_��Q��r~�	�qq[����F4��Q\��ص���ke�������Ҳ!��d�6�:���1kݶu�X1�1����m�v�X��(Q��\U�p���������+Q3���y[�[V�>^HLז�.͛���֚�r�<E�F���i�=v�B|�5��k"���w�����L���Y�ؒ�z��3�{ ^��.��k(S�9O����6�S�([��,�`�]��wN�%����H>�?����|�r����6�L�R4��_h�Ҁ�DG����ǖ���C/�B��j���!���󹓓�r��/&���g�V��e@Ơ\۝�߭�{��Q���=�� �
fo�6��VL�)����K
�WU�-�d���Z��z짶���A'�-���im�#N�h��ݛl�49�`[�����0��=i2
���8z�pk����"�U%�#�d��������5��b�3�@9�V���Bm���N�e���Ύ�'ۣ�1-��=�����l��	�5�;�$5��=���c\�BSH;2�v�1&D-sz�:!Y�]�m�+)ϡ��O���ʚ�w�R����'S�U���~�sh#oߠ6�;7`����ߗ2ͤ<^8����t��H�lL��M�=�����+g���({{�ܱ�k}��3��!ʹ�΁k5�~a4}��!��₭�	d�^�_��:ў�n�$���!j�Y��#��8W��/y=��HKK;��%R�KC�]s��R��C�\�.��9�ݢ���te|/��J���=���8[ xff���X1
7_X�EL:kQ�]#$xS`�l[j�M������*べ��u�������ܱ����;&���lgV���**'C�S�_�O{~�@}eP�3QU]}6�]��v�����ѽ�I��]Z�<�'ݨ<@�`tD��KJ],�̩EO��mʕ_H�D��1U��?NG�hM]�ϱ��\�iK�Z�k��ы�ł�'�W7Co���:�`O�Ng0vvu���Zym��^�;;9U:�d�.V}�H��������d�%Q�����/�ɚX/��Y��8�W{�@�s]�K��5�8��!z���r!]	^w򍍤�Wv����O�a�������<�$�8\�=66�r�Ն�iwW`�fi��v�^�/�����iY�Js�X[g�8�������S����j�Vs�������������h(�^�Q@g/oР���e��� }=��X���й�a=���p-K�����l�z�F)��T�4?ĲdX��O��<k�r�J��>�7����o�=���0���P������J��ö�]j��?C�lM�̩�6��u�PҚR딗��d�n�91���
��eϮ���t-��?R3�S��4����G�YTm8c�N�[�)J�ν������#U�uuuМ|�guqE����b$�-	4����9�jJ2V��Crn���f4+6��>��GP`jjj��õU��?�_�h�>��㙪��k�F���p9�:�����_�ɘ���P�Q�Z��yP���N�S�hjc�ۋM^��t����맇��ˋ�/�,��c��y�,���s6��lv�9����tS�����
`e�]��(]�P����QQlH��� �U/}6ܘ�h��R�9mĘ�d��f�$���4�[i_�]_��)�tw��)��������/x%�߅��T*_O�b�V���}J�س�j@9��1�����#�2��μ��sԎ�l��4��TR �~j5hju�d���|��O4�\`�4���W����0P333#��J���eftv꽯7a�C�&4������@�QhR�6Bj2�~R�i%.&����m�p��N[��[���.���u���� p��sSRO��	`Z]�������tG�?i�����>H&zTKxn���p6(!o�_u��d���:��3���5~ȕ���P��d�i �2d�k8�~Q\]/;���iy��D��_]]��g����� ��ۗ������f���<q8��?�j^'{wgN}}#T���	4s�sV_�\�{Rô$�4Q��{���~�q=�mJ(QU��-���7>�p�a�jUԅ�Zf9=j\؟^ϻ�sK�Q�"f�\k�[���_����ƍV�L������J]G.q(ΰc�^��b�@��D�|�׹\�ܭlI剉�@!��a���gΜ��033�sT�*�� ~/�2�ATWww��pCn.�����yc�����������Y:��glH ��+*)�?{v���,�R,���L&���H�3�b�^l����zzzofX-X�̡�4��dB��v<3���(�>=5777��i��-X��ǂ�%��� �0�2c0|�~Sߓ�t����O�r����ϓ/�Fd��K�`�c��s���z@B?��z����($�A��x#G��nF�:d.� �b��J����V<��Hv&����lgCj�i`���Q˻�űB�m�#Ma��r�TjKu�\�ˍ^��s�$+�Z�A�	��ŕ�/,��1�*��xM9M��G�d��d�A�W,�5�M*��þt������8�\�З'�ي�;׶�|�������(��� tv��ܼ�����&-��?��?5��LWW��/eۮ��/�er�G�:��:- %��y/�<Ew?��j�R����ِWZZ����K��}����ǳGmI�VZ[[�Ԋ~����^=�?��Q'���={����q��{��@����su�N�]����h�$������{N�-��'R����[��ͱ'��q��<Q����Q�B���A��%����n%u��z����͹�v���\~�&ό��o���j���gS`)-��"��	�����9b>�
�OX/�Rh�UBq���3}��J'�����0���'�*  ����^��b/rC���;��/n�L��S�cf`=��Ҍ�-�M�nħ֦�~�c���O��Q }�����H����e(��q	�x��E"��R�|�
᭫���:���߫s�\���y9������(�]��*�S�+=�9�N��瀱��������a�I��{�6~�Ħ�-��Qi���� ��&8���db���p�唕�?~� =ǹ�����Z+/$�O}ȳOT�� yDvnI�Q�X���Yu
f�]���V�5^A5@�u�Β��-3Ù'��@� q�T��g";;� `���v��b��Uy�����.�H,7�ua�[�4��ұ�þ�$��ϋ�a`��P����j�q���[
=#�L��3YJ5Ⱦ(����o���{�x���}�Q��;�Z�K������/ġV�ΥБ���phMΞ�q4�ąTbk����ƛZ�M�� p� ���wOO�l|��ZM�B��!�%ڷ�=�Ll~���5 ��� ��3h߸�֗�h<� ����鹨Cj�t}/zf���̀t4#~���P�!UB�X��6	��K����=���&��,�v���-;�e	�r
��uF�e����`�|���o�O�����P�9�6�W�RI��Q_�m���C�:
�������2ٶ��Z�U��S��\SR��#<L�EJ��y�yM�蟹�}��M�{�4i�2�>�|V4��].�B�y˜[e����"t�q�_W|ȅ!u�U���8��Lmm%55)�_���������Q�D^ޟK��T!���8Y5�����@6����
=���g'�{W57��5U��vil|{��-����/~ �&��⁢Ǐ_��>��T=�����Z"����5��#��>���o�1�J�[Q���|7n��>N�_�	�f�]�Zm��� .�'�$`����!X�Q ���n��5���X�t�z4T?"�T���,��2$��K@g^������h
���X ���r����a�aLH�e��АÓ��p�r�8�rnccc�u$Z9��$�Ӕu؄7� vf``xY+����a��[?��ɇ�V��� `�$a��ڀ�{({�b�����UFɔ����І��Ng����������[)�p;"����ҷkg���|�slM���-�!�a]e��>>�@!��mU�^���0�+�Qs h`����X�J<��c�0�}�]^.@���tfSvi��j���/�Å�[7u�;�GB�WM^@ɿ��Z)8<�7�r�5��8�����,s5��ҷ��,���M�@����;�œt�:���Ҳ�����pN�tT&�}�~mt�(X?[������j�¤k��M���#����+�^~�F\i�]eGj���ߙ�,j�8�|ȍ �իW������d_(q��xω�@���F�~]�^L��������{MK���><-�&�4��4��K�苖٢QQ8���%�cOJ0C��g�12r58����텇��,�pa�o#��絛lJ"�n�>�tF� ����JS>��O�@�2Ny#=�׮#�!�y2eM~�(�,*(�x�?�uU+�=\�������Fȥ;8�{�ahO�'��痖,""�O��Q���'�T �E����h@�^����p5��H&�TV�q�r���\MG�y4w��V�R[�=�b��a�I����qC�U������lH���}�|!�뒂Z�t�6�Ԑ�U�_̢cZ� �����S;�n��.����j�CVҚ'"̊�1RHT�b��죄����Zs��س�I:�R�%U�%�E��섄���)p�;v���g�H��������2��Ѵ�Q��� ߛHUn����@|��(��6�C�Er�^/_uQ`C�7��Y&0p�_��p���P��*dR���u���!>�^������	��k�,�^yM0QΦ��RCbЩۉ:?��6g�Nܱ��򍃜��_�Ϭ���[�93lcE���%^����	�܊�S�ڗ���Ԓ��#-�dX.�j��ȡ8״M�Pj�{��� 9����YYZ:��t����5m���7�&B�B���ˠګ���y�ܚ���*~1�O���j�`*�F��Onz�,sZ
�%A9V�6�,�E�+~��#`�r�6a){�������^,���
(K���f�~���. \���,��ڼUUgۚW8O�z�?���X$�c�B7?~� >��e�5Q�驏yB��Df��I�<�KĎC^��.n�C[�U�xC���g��l�`϶����a��{k@t�	Fxxd��_��h���u�
v���rHc(��z��̣���4����Vm��E�մR�B�02�s
֣�߰��C�lWn�\�S���#H��s�{�>�M6(�B Y8�;�y�>e#�>}��l�(�v��	`�g�%1�y�Kp�T����<Û#'���A���a�!�7~M���o�zj`mt������+t�����X/̞�x��%_Dkjqkj=�y�IJ�Λ�+ŭ���u^�5Slp��mwww�����{�](��G�wG5�m_QP�*
*M�WA�tD)�"�z��Wi��@��Co�ti�w�Z���x�{���;#��:��{���<g��.�H��7���Ձ�'�㇛^G&v�G�z��mV�u���X�A�C>sraX$����f��"*Ɍ/@N�8+����3i�Z}� w�j����g�m����$��;�Ȋ�i�	���˂��l��:�y����0S5��ͅ�Ψx�D��-99y ���M/.5
&H+mDx���y �@^?J � H�p��٩��1�tM5�9�����>�/W\�0���t�ޣ���vu j����>��8$K���A�%�DtC=�&�>Ѡ�?ծ?d=�o��W<_	�P�5!� /����̄�����Q�A� ��ҶṺ�����k�U%L�=$�g1��؏>ܨu���M�}��@�y��
Xxtm#�s=�H�!���&~�r1��=mξ�)S�ֺ��H��a����/�dn*����x����GL6޲X&��ȪC�f��j6p�����FjD�ڜ'�t��S��JJ��O�`_i�kul���5\u&{u���Qo����1Rg�0mVO�� F�sO��6��WQ�jW�^c[(Y�6˱4!����̺�}���WkNM(�
^���<x� �q�$1`��@�;��d��8�.E��;[���t��7:��*��'��#vD+�XEE���u���o�ݲ]��H���'%x�:$�p�m�06��gYh�o����y�Ԫ��Ґ��(]�΄�.gܖ;������ׅ��zd����]�!�`hr2����}˒0X����cڠ>(����U������0������8����%%gr7'CT�� D�:�M`�n���B���W%>��SM�Z��"�[8����Ĭ�ri�ٴo�����^�a�}Խ�*лt�`ƕ���m.:S@��(>*�D!�/�\��ƻ��TB�oo\��^���/�*��Č�2��´_0�����#��&�rUm�r=�X�mOZ��.�a�G���:��Q��Z��獰����6��Q�d�鱩��:��&�Ǐ���WH�~�-�r�z��H�%�&g��5����Tݒ�����*��c����缐z܀Mn����r�@@xʗ�d��2<.r��9˱������mf�!�Ɂx��]��͈s�9�0�]1��"� d0aL�k
&���J��(�U�H `����K���g�� 0j��jmm��~9��t�]�~���a3~&0p�N���o#��P/��H|��4��O��tu�,G�X�����R�PC��i1��p��4"�3��$%�CC,��ׯ�]�s��������C���-�PC��Nn�#ڻ��%�Y��7�.�M��:A���sċ-�>}�/���T_�u���k"�C�<�g\o������ram��5��C�/����o�Ex�nkhh�|�:02�[:ܠ����uh1Wo�b��j�� ׬1bn� p�F �B)h.T�܉�xA�@@,aA?2�Nw�5�%���^�>N�`����8Ghh�j�� ��!�]`�(S�3S9���w�׏����fq�R"�)�:�_	##o?�ց��mYI�1��Lr���0ĬH����	+]��0���O�H�&�~���H��ӻ�}��y!�����@W�������ۿ�ۜk����ȑ����yyK�,�U�;�Z�2��/d�)�$#0���@�X��Je^lF�d���� ��z�.� p,-��D�����e����Y$�6 ހ��w'��A����ېSYY�05LE/����u�.��_�|�~�������0)�N2����RB�"���Xw1q�Sօ��=i��K�3O�JlQ�S��)��-셓���3Ņ2#�;�=@~�R�2��{�qVL}Οh�8��ɿlW���h\�5���["��=x���zl|�9%$56:��d�@�Y�	bl��� y�Z��1����>�[q�����~~���#U�+Z�K�:�:B���TI_���1��rRz� �d<,"�#��ҟ�8A���x� ��J��m�	�� ��k6�2V����D%6!�?p��8�����G4�-]1gC]q��0Pޠ���Kݵ�f-���0�a^2� ��5��v�H�
��Z�n���g�֎�)���/W�h�n#� A:�Q�7���p%wO��i�i��W�e�'��w	s������^#�������hL9`��W�>a�!%~n���_���N���'���k_�C� �P��[G{I������`OU���� ����0�W�*�v�Oy�m�.�.�����$�����A�փ���t�m��ʣ+Cx�%���H�M����Y;���Y{o��������?�����jJ-��U���M)�^��,�n����܄<��FH@��������|�Zr����?�����1�Cx\0l��[� ߸Tݯ�������U!����kxnz-�%V)'V5/�)k��;X�� �ѵ���~�Bj�h�5�F�D�'AE./[g��&�5��@ٍH���D��{N{��`�����"Z�Z�i���h>��	��ar��������f�Cg��Cɉ4�r6D�S.��������i�H�'�o��q�B�D���^����1=;��`,Zjb��(P1��Δ
��w���A�*�����)�i�}O!@mJj�uU�3�у ���O ]]�d�:ұ�~_��Q��Чť%!�#)o�hE�ħ���M�D*�M)����o�~�z��y�P7ˮ�a-�ccЕ����P:|u�B�/~'��|��ˉ.��a�6E�r��::��Smdr��N��ۻ$��?b\p���Kx�LY���H��}Eհ��gFq��9�t�H�È�U��>�C�90�P�&���ob�`�cE�����r������4S�����c�*���l������#�=�=���n]Ā�JO�<���h;b^K4��M��n���E�~�JK�;rr�[bd��Z�I*�:�@59s�iH04���#�_�?t
�����_E_9F��q^W�����ǫF=bcW�Фl��/(Z[/��Z?��Xf^��Dc�g�Z�l�ix��3��L97_^Y[R���٨h<�����SO=���C��[�~WG`��<����6K��tP%ǁ�ʻ�⦧���f)�:&�p�%�1'��� ���А@y�3( 4��1qj�~�\�6kP\�¼c�\���@^A���̃�B�x�I`XbI|Z1�ڴsaK�ƭ�#F�;�7� ���{�_�A�:zR�	�ql Sn��+[�%F��c)��,ĉ�"�I��ib�5�QHz@�^�����O����Ǹ�h��l�=�&�|#�#ZQm��a?�b���ǽ[���h����[f (t�2�P���`��Ʋ�:jH�6�-���?�T�/Xr�9:�51������ˤzڂ7-@���K�䮑,p���"ZP_1�5L~qt�v�~�`��A�ݘ�U0�bg��g��@��}(AQ6 �uz���x�ϩ�)�leK$��^.'��h������%��Ռ��1C	����X�	4����I�B�=�߯/tm�"���P6��wy�Y��բ�D��5H�JLLLZ�o���hUa���&�
��3���Đ�W�o�h�+�G����n��)-8���@��-��7T���y Y_h��w�{��~O�QdpB��S�+Y�آ^??���h6�p�D*]J ~�Do��CgѠM�8µ�����!�=��ߠ����f�x���e{�"$���צ�ѷ��S��r�_Lv"��%�+�7;�oh�m��t�xc�ֽo� ���� |�����@6�K*����hi��m<๧�?���^I�^�j�����v'Hfm���D����Nfff��(�/ο�@`-hN�_�N��F�(�&�/W��p^E1�pQVL>��DT�� R;O)�P�x��
A��'��BD D�O��g+�v��DFxu�"+�?EG���C�4~���BXa!�e*�C{�TU_���&^i,v}�8Bg�4"�U~�<�ژ�J}OKpWB�<&il�8�h8�ڮȚ��jNd�������U�~��1E�3a&$F�"᪭���19�"M�3��	3���+.��ц���옗v	�c3�*<��U�����{���#�jL��%�%�C6�����6��j��+D�2a�}T#-�]-dj1M����Y|�����!�zkfڄlҩ�����bNB����Iָ.��Z��ۮ��<����d�]�1�/��ȯn�C����6���kʋ��|�\RNlQ>�H��W���0�B$����8I�O�w=:�!C���S��#0�j����w<!vހ/��ob/zxgb6��<��L4=a0;�8��|뢙�7h�ǖv�þ~��sO,*_�l`�ZiMI>C�^V<Zb�HI	�{J���uR�o��� lJ��bTN��������C��YZB
/��'L��o��� (K�1Q����'|FE)�|38l8PHj|x�8$.Ņ1~�H�#��x_��o��7����n?�oS�����_�����4,ͼ�&'5mC��j��I�ג��8k��C
 �4�K�I�+*�Q@b�͑�<�%���0JlS6�/~#�g`׵ ($$Cm�]/������aC�,���\zt�(�>*5�
>��|P�H� }?�A4F�;,S��T�p��շ��r̵����U��ۉ��n��dg?���K��@F<i�'	cdt��q2 ���H8Q�K�lF��~���Z�A�a����[��<���lZ�՟*�;]�;���
���̩��+:��ɮ�)������h�/R�?���po<T6H��܎j+�Sb9D��p�z �r\� <$F.�C90��f��}�A*�G�Y��ܘx�H�V�8%o#u��~I��ΗeiQ$L>˳�L�<����")U�ٹol��D � >�~+�;���2�\ ��܄��7x.3�sF�@�6'����Ջ�'�een���Q�ɩ���Lo�*#���C��a�ÍZ��M�!��+����<��D�֣� Ji���|�x�]г����Ӵ����GF\ٮ��g�7Գ\/������Ѧ�<�ĕ,�T
�7
2�+���j���r�!?����A�a�Ļ��Ff��!]�y[$�_@Uv���󒏄W��dhi-^ B�Е�j�X�����p���˲�ϩV(g�{��r�������ld���p3�l�C��R3�h�&�5���u�L���K��Z�Y�w����k�$D���F:���1R��-W ��tFCC�]�7Q��: [�]��^�])?�߀<6>ؕ4[��R��:`D��� �w��}r��T�g�)�{9�6tB�M�9���b�!Կc��<G����@7��*<��\0��9��u�P�?v)�;p*`M|���+������4P��'�����O��6A�7A����<& ��l /�PSg���:͋q��T"f�dvZ�7�^<�f�B�}��N�h��-���&W@Bn���,?<G�T����f���N�i<ف7��%t�o�n)c��G�aVYW�P#:�j<	]Jy��F�Z=� �M��� ���ݨ1Q�`0�1�i��"\\*ܙIR���M�^�HJI$(B�f¨����"�)�S����E�O� ���8�բ
q��  ��t�ˊ��;b��G f����	���2
�O�`�X�s3тt�r2�.�֢G�ՏZ66@UVMU��%��\-�+���&,��![�b�vll��k�r��25���:{�芥�Bv�y��w ��M�y����^�]���4@}���#/��d vO�Ӑmྲྀ7����nnn���^?�g��d7 �����������7��s1�B}b��Ș���i6LB
j�C�� ��1�f��")�F�9T���1ZG�K�ٝ�b�t��������H}��cz��
{�d��f�{�%Ȇ���,�%����ᅊ>���.��� �ʹ,Ɵ�{��f!9O��]����pD\~1�#�q�hG�� ���>)1X�p� =�C�3����L].2�d�b����{�+�w ��m�"��/3��Q�������p���"�n�{�Q��w�s]�����DK/�Fb��B����)�b�p~�W�ϳ?��=.�����$r)�3p���q0ρ��H�O���.��lDmy���1}�)7B6D�R^�=7�G��s ƫH�&i�&x�0���Jv���y��[���E���2mT�F�i������gpY7���Y�C3=U�3��|3�%&:�v�ڪ'�7�STڑPi��ũ� �d~�-�=��[D/� �n�-���:��ބG!�\~��
���#��w���堁<ؗx�sa �-⓳�&q�X[ԭwI���@Ä���ld1�� !���dr4.�ԏiD[ ��)��g�Si_<=ۈ~��i�Zb�q�Ч��I���B<o��9�4d�Ү<%�M4Oi}���̞L1���ڑ�"���R�K�W�}\�yt����c���'Rw�t��<�Ҷ�M���zr��SSW��@Lj�8Y(֝����)���o�N�>��s��BH=˩-�o�L6$�+w߯�獴��٩�$j�~�!c��2��`���?��V�0�*"�'��� ��<s��U%�2��b�2
�AZ�Ԛ9�]2��eh+Y��f��)P�UZ������HHS��Vcv��8���� Oz�J�)��h�����-=ν�����nB.ń	����\�@=ٯQX����!��eL�iJp��;M�$$$�猛
���d� ��oȭ�^�h9>Wf�ۡl����L5�ݏG�)�25#�q�C�6��+��f#u��-�K?�(i��(���گǹ�Y?7O�q?���~�L�x��aw�	��dc�?@a0��C7VSs�F!�w1�����Zm%IH1k7���k��♏L[�؞\o{�Ԧ�Sџ��(�~���ȟ#:o���Xʭɛ�FO"��ҥK�?�0z��}\Q�����-�U!�����+?O����O�#f�9�Nȩ�"�pYcK�)p��c"��q�G	��tP8+++%w��p���s����@�X[[+5\��z9���*z��P6c�;-OPE���9�N�����d��H����>�����˝\Eu������ +��1�6�멹D7�O�@�BM߻�"�U��}����=g�/�ꛨII��gAg�s�h��ʼ��X�([ *��ny����f�U��Ǽ/�r+���2��_��2{n��!�=!��3�.��31{U�����sz�����'�����2\����$Mv���M��$��-�ꀿ��-�|F���D�)��V��X&��A��?�0K>B+0KrcH�=.����oX�B�ܟf���:�E�����1j��'�<uD:�^���P	�+��.����G�?񳶠R�A�րD
&�6�a�>]���Gd<iry��U2�ʻ��u}A}�fȵV��!׆so�@T|���n|]��)���lFkk�Q�����B��
E�ǫ��w�g������R=ryt�����ޱ� �I��ы�ܧ�C]�0�5n��:�f݊Y���mǾ��}ll4��- ��{9��ѓ��Ӗ�F�u�`���d��1 6d��
� �ۄӼ���g����e7��Rm74�F�.A��&p�U$�9����g-x�(�w&���N�E����`�TG{������x_��"���p0��]���G�r�D�ݵ�p�>y���A�om���s�N�[ԊX'\i�\?rTS�կv�2H@�X��.�f���k�����#�l�3������^
%	���E�����>�D��Sr�F��g��� ,����(��������O�"K�A�ӵ�V@�>Cں���?�-��Q�'!;��@���#��5:hM��	�}��g��,'Jd~��c�������_
tC&�.'�)���	�����e33JJ�G�㍏�_r��;��p�]c�?e{m3 JS �p����D���J� a��@�_3F֢��6v�6��������Ϝ >%桫�U�xKe�#G�V;ٯ�b�I<k�D7}qz��q��sj%���������X�+W�dH޻��Μ{� hɍ^��0�R�1[U�ͧ��q�P���'���b`��3>g͂�z�oɓx{�E}}�Ҁ�;}�[�.j9��}�km����w�f���&6�����V's�G]�xP��D���<\��o;U��]��!9����Lv��v����[e�+�o4���}�!�S�\��lE����g(�d
6%�?~,��+C)���'��-��󵩮��]Ko3�A���S��DT��Q������bѦ�"2�	wO��ē��a,���3a�#f�)J9���&�����A�f��΅�ׯ_�?'X"�bxB�K���y�Z�7PnK��5����+s1Y��X]���{)`�<^'0�qp/��_0r����=�(�V���ݟ�i��q=���7(I��c����pw-ޠ3�k�v����>~� s�d�BNT�K���4�{=#�3E���TWdP�)^�w��w[�C��K��X���I|�;�Aҭ@O�X~��vݿ��r���s�6bR�]�a��F���:�#&X�'����qG�RXҬ#Rr1��Q���(he�));i�5��q�kޖ�R���h����[A�]���� ~jqڸ���Z|5#�[?T�HO3w*�l�V��6By���3�)o:[BW�om俼ə�܄�	�U&�j%J��.�bTg��un���R2�=��۷oY���l:��[R�Eﮍ=�ä�u���96!�}��(��}q^����{�k�{ON��b,�&-wl���7���e����{���y��D*��x����M���V�լ�F�5H�Q(�����"�V�����T3�"[!)W�ZZ���K�G�D���@��~�B�n��T6��CRR���p�ѡ(����(|���/pa^��0e���mxEo4�H��j������Y���+g�ҼId������Q�����,��W���9S�,��-��g�3�T��J�)��*]}����!Apq�s����Ϳ�c���Z�|)�|i�(����&:�s�,��²�7J=��eW���ݎ����}��߱W�6�����A �&h�6����X�!*<l��.�'�S>���rc��܏�lB��IO�=����D����a<�z@������ӑ��&�H+@�ThӇ���[&�RD�8J}$YG�<Оy~������=��J��/��qy�q���J���6]}#�u1�|�$�T���	5�'&ބ�`<ˊ��Mx���ڜ�G�!�T	,�����O$���7�1hΐ�_��T��*=a9���+x�� �2vȈ~����Z�Rut�8��B���E������'��}lP�N懺S��G�؎pL�;�u�Ol|�����A��7���v	hh��(]��c`�	6$����9���%NjrU7���B^��7OU~��qN�'hOftƀ�̪>����]h�N�;�6���F<�e�rf��*���0ʌfh)�w�R\�¢RH�$�q.�Qʸ!-'�|z{(��3���6A���F��'��Oz���z)5���K � '�YJ-��;8\U$`�?��Ml����ZR�K�<}D MN�i(lxX�`S�y��`�`̀���Qu;�f�i<��Z�H������~7"<|r���]�3�E#�}TK�`��[��⁷pt��4�b��i�H��.q�����(Qڥ�0 ��r��1��C�����:Gf�'������S����R��O13e�/Hf�����+��/u�G�%8��xυ27f�@�tmrU�7{Xh!��0�,T������<��Vǅ�����Ȏ\(�zC���`e�y�O|���V�矶)ڲ3ߵ�k�Kwؾ`T�/�#��H��}�3����� �F�0x�>�:Ǚ�u}x�G-nM�Y�8G���c���|@�D#�In�/�zT/�*�R�DW��:'�_9�fڗ"d{?�n�S��tݟ�-=�R��������J����(T�aL�q<��r�� ��`*.�b��(F�-Ne�������Z�~������)���T���_&��i]�ϔ]��t� ���]�(
�����Ng�S��<f�Ԗˉ��o�̊�<�����T���rd������>���|��4ہ)l,�1T:��P2d�Lp�}8̧���'�)��Dm����`a�m�s=?N`;��V?��tCSE`=��K��2��Z�-\/�`�GZZX��U�{��%4���Mx75���G���eB��_���a�Ӎ"*ė�,�MR9�{�=�ɇ�_�f�����=��� ��p�?�s䨇}���׬�\��Q]Bm���A���J�W�c	�(��p��wa�Ú�8�-�L�bצC��W�\^�
ag�ߋ]���ͽ�D\�[��{���#���o�ǩC����7�8�tN��k*k/ m�d�H��dPs�*mH�B�H�6�χ�߯�uK�=��Xiz[��c-�6-���o�O���n�G�E����Pl���؅ �f���c��<|/��Ҥ�=��&;��͆����yl<j�뽵�������۵3���{B�03#���3��h�rhĵ=HA��f��)n�޻���b�uo2._���n>�_�5H�QW��C4v՚�8U�wQ/�9EΫA�_2Gsd��~l�_a V}%���8���#w����@t3�^��7�]%�5;�H^�b��3����'�y`~>s�l��FF���#�HǑ'F���p;��5c��o*�1Psˊ|� ͅ� �+c��'�@EtØ%�n��Y_�ڭ�Eaa�R!]��Y72�/ad��aέֺI��1��T�����o��^�i���x�%BY�s4��b�*�q�*$��A����jQ�|�;����'�0V~�!:��s�����)4Y��հ�6�Kgv5��_����c2N�WW�c���S7�d���}񹔆��\M��*�I�Zq�w8%�=&iߧ�?�&�w`��R�e���XA�|Sx������|�]c]o|��/�.��ϜP��ߢП�gԌ��~�m�=��߶�R��]���ӟ���"��x�:��|<����'iy�(48������]��������7��&����
�AbUX1��Y`�=���!�^3�v]�SB�?bD(�&a(�uf!���Vc�+j��a3�H5���U	P��l�p��7�'���|VXHڃc._ׄT��_;y��	��[�%�c-
�}Hۈ	�/HwN%d%�N���0�q�`�y��NK%�e��v����N���<{�����#2q�?�-Fsb@U��(�#�@����}���l����ۜ�n�O�	x*���%yfk�֬�Z���Ϩ�� �*78�Îb�<Z��i_Ȩ��h������k���8�Fq��3`��=Y���p�����R0��갚�ḃy
�ˌ�]W�UT��'!�F$�.��.�!D��U�9.��R�@ڗ����|��
�|����Ӽ��_�>��{_6�nk���j���	�����:A�1���N��_ nK��=����9y����F`;�^`��Ⴔ�B���L�o���՗�4�$�O�s@q�뒵���ꍂZ�%±�0���K) t��WY���R�F��'����������,�t�f�gL��}ڬ��6�6�Є�)��E��
��U�6�8WE�}���au�����y��fMě�l4����/ƙ���QZ??QD��, 
���]���{�L�q�����>?���4v9X�ɝ9������SK��+n�x�a
�d�嫯)�`�r��4�2����˶�ҙ�@R�J����:���������~Bk��(��<��洮����ɯq7�%�vR	�3K4E�c��N��؃�<�U�!�=��M�/���U>9��w���:�|_瑟Y�J�y��l��pw�x���ȓw�M��&�q�~�k�B�����Z�^�m�T�3K�*2H���Z��N�9��u�;a0YN���8���s�s��¢n��J�ez4>}�q��ٿ9*N�xP���*��s�{wAe�byܾt��w��r�bk;m�G����wZ����/���Ο��R�_8x�V��V�q��Z|�N�K���=U�����/�S�oWEF�'"�X������̞Lw��|*ӥ)u�/2+Fq�ǫ!��}�ǽ�z�]�c��AU˺qK����ɒ��3ݱ��нR�u�}�π�7/���]���d�mՁq�c��-��=k��J�٫�5h� ���Y��r$TM+헿ךlƨ��=:����=U�"�n��Pem�p�
1B~�x#��Ke29齙�'��~�H,�V�Ԉ�m�D�	��e�_���Q��5��)�%���;�0�� (��d+����줯�K4E�0��S)�Ǜ���Sw��h����PoI�v��2��#{oI�ԫ���*�;����mh,'�;�S�n�F���lM����՝�ӖC�pVpPj}/Ų���$|a��(}C/'B�؈��OH�jﺾJ������G=0�3��Q��$�zz�]��,nN���R��f�Og������DLC�a��A�ԓ��̡�aȡ��&]����C�� R�����}^��#�����Vg��~Tw��W__K�V�`'�?�>�*r�%���n�M<���p[$��w2?`�7E�zb��`�|�������5P�	��l���bu׷A9���/�$�?cʡ�u�^(~%m-o��6��������%Ѫ�8F$p��*$�|18)h�_�g�Jav��C�Vi~J.vR��7f*_�G�su��ڻ`����s��/��
�|1���*���Q���@�k�T؍��TW�p�W��g����?mP>�`z�y�Gڐ@B�_巣`4���Qۃ�Z�;�-:�1/z1��p�S����JPK%�$�!�������������>���M�W �F߸�����ӡYS���%���":7]�~���>�f찥��3D,����ٰ,p�,@s��`��_/�Vc��%����U��a���Bs��Էa�r�d�c��絭�#�F��L�ۧ��G�2F���
-� u�}a��<�P|g,|AH�!�Ɣij���6��ĉ��V$��]��<6�.7 *��N>��k[�c5,"�u�n`��<5�!5�o�����<d���z�R����P|��8�Ɲ�0���N��$��Q>��z�&.�o/߈�Rئ�'�d,�u�>H+���бƮ$�����^>cC�m̔k��p������U-�,x�L��b��q���o�A?g�������юh���,=3�'`��<��O�ϝ+E��J�,�+[{|�������V��xNF����Gm@����`u�X��o�)�m�����&�P_�,���`�9/C�=�g|ݸN^C�������*�-9.,9$��,������W��OE0Vc��n��k��4 �ԓ/��	&��X,�W�*�r���뻗8�oYG랉A��UBB��V-�#����˜��S_Ɠ��oS�)AH'���Ig�b���O�������`�l���;r�7Ի�:����m�m�:V�jQ@"�ٌ���j��UJ?>n<\Q�wy�X9�|�&��)4�!��2!mw����fO�G��}�����UC��Coķh��Q�mhj���[��s��)`��N�tӗż� �s��OFE�9p�:(�������l_{=�F�?{���_�<�s=s����j��&���R,�#��s��6�ثAM�FEk���"(��*p�p�1��~0�7+d\a���u���������p���*kڂ(5��m��J�3�#"~��?~o�k���ŹXP�Kŀ�Vc���V�fm@���'���Մ�u�@LK��R>�XԻ<*�$Zm��pX�5T��ߢ'm��y��w�B�1�k��²��⓲�ǯE$DN�f���7K
˸���{[/���6�ɝ�����om5��6tⵌ�Dm��*'�K�ޮ���jA�0�P�Ju7�,��;Nq����P�a7,��ȖA�Oٻ�啘�i�32.�����;z��E1U���]X	��������0~7u��N��2�*��{���A1�?o7d���z������v�/�;�h+���-DՌ�"�ޡ�\IG�Ϙ�)�O�j�U7<�j��@K�R!������T'�R�-�������X%�D��][�����ӭX�T4��Y�/�M误u䏓Q�>o^�U��X��vS��h��~���I�`Rt�w�g�͈���Y�����/#�3ƿ��wMx�1Z�����nCF�U�9p	k�=���Zc�Qܺ���ZtR��v�:}Cl��d��4��^_]�Ή����D��2��?s*���֭�Q��9{;l(R��Y�����#L~��P�\��1���%}���c��+�c;:	����/�vm�<d|vC�(O�8�t��˪�&���!���(��B���>�"���;$8흩X��Ŕh�缉޳�C�;�Y�g�p�D���G��V�������O�uy嘘�:,i�׼�䓊�bAz��6�ڿ;84����6�=�*��D>~�c��d&��p�.��P��a���r�U�!~�eͫOi���5Kb������CY0P+�[I��B������_=�U���*i��o�|�pV$���º�L�b5)�Z8Q�4�Vu�z�f�8]u�*�q\JP��J�*�}�0�\K�O0�~��P�����O �qY����o�W+��i_�ܜ���:{ ��mүуL�P�Tx�>�]�0�s�Uf�P9��;�����=��SS�|����r�Λ_�&����&�۞�]�]�l���,�z��C��ɒ��� �͐g��C[_����X��{�J���k��rwN�&�6ė	*��n��A"J�Z#��os7���jy���\�t�:�c��_d���U�-���Qo��fjLP����U�XA4+[�q�Y��b~�����qa��'2h�Ġ�ܻg�e���lY=EA�2����F-{�lZ��l���������w�_R�1�3��>%!�6SE�"��ƹ1���ua�>�xːü�_�3�-;��s%4w͑��1������P�n�}�CJ#~�1���R�E�;�>5Ξ�n}��q��"eK˄�eF�͛�Q~���bU�^���/�:ho�u�p|�w��zk�E���q�a'qO���ɬIcnQ?����"��q]3��R�)l�U�׈%�hD�����V��L�z5�ŧ� ����WC�pZN�gN�М�g���R��ɭ(Y��ΗP�_Z\%.�|"ehV�ST�t8׭��5���~��\��GI�����:�_���Lk'�-�LP>z\ɖ�9ob�D`��/ף2�T��9�:�h�=��ـp���e�z�n������h�T�G��T6�q�̞HY@���jo\���}�����Cv��d�x�.�d%1��S/OK54�$�����G��3�\����.x��y��ͽA�Y��w ��ֲ��US.�D��s�f�?���X�;=����o�0��	��׈&��F�����N�T����@�2�NRt����͡����/)��9s�
��&��Q�u�ǽ��(��l�8��t|��k7��������]��_���ؚɂ%�b/�z?�x���5�'9ƞ��w�N��6n֬;�FZ�Dd��\,�)���ʠeP�O�����^%��SCbڜZ�`m~���r\Q�(.��l`�b�91�8���P<$%q*fz����G���>��QB�*D^q,�M��<�$~���ɇ��R�D&��t_�ת l�2�����mQT)ۅ�u�K�e`AUtQ��б�χ�M���wR<}������u�tZ�[+��
��s�JJ��D"�r�?�0s��{�>^�/���|���,^��(�{y�?���F�H�M������I!���������\�i�h����*��;����N���(Rk�'��a��_��0ń�Ft��t|�8��gz�V)����(�aa^3��mt�L�����]��B��U?1�-���#��%�PoY}�{��6�cOQ�/�41�f�Ǧ�ecg��l�>2j�Z;i?��WqǓx���'ٵL<� �U�e+�1J�K�T���R�;D�Ƞ)-��wF�Z+U\,eMd֏4�_8MV�)o��o�m��� |��!2��ߒ)C;eP�®�k�[m,�T�)3�V�6�?>�y6�3vA���;���܅�ѥ��*�8�^�5V���{�;��K�	zП�n��u��y025���/V6HvƿQYu�����C弟�`N����1K������,I<9���|�z�����w�a�(1�ŭ���vy�d����]o�'R�`�k]X%V��%�JQgn	�#��U����N�l�����ܢ�ء�<�JfE����,��L��"�h�EW��@���9�pNe�.Z�j65�ٖ����:�I�R�����b�ȱ�����[���O�ڤ��y�L���E�~���,�h�N�N���PR�{��Ĉ�`������Y���7��qUV��{w
b~jr�
���u��-�i�:�9d�.)��+����eۈNt���Vqvtnw��V�3F�u�=m`N���Z#��|�7\�[��`�X>͇yWMl��0V�9l����t�M�g�r��ʨ��O���0'�)W�j��v��\��M���V�/�(��<ȃ$M�Мq�ʥr�%�U'�s@�%��ѣ݀�elˏn��,9.V7�z�S~L*��O�_ �N׌vo^+5Aw1�k���#yS���wh6���	�9_�ԕ\�u�$��o 7��I5���GQ����+ 9�QrO��ڟ	hH�}��/��\��x��2o�� ��i	��j?d�u���X��%!ɚ��c�p���>s���En�0��$8N�=�M��k�[��T��>�쥈��×
��m]�)~�H��ȑ�~�b1O��:˱�����>X��8����������lf ���{ϰ(� \E�EPTT�
"�!LdQ���$�!��dA@�"   9*I�HF���3[���{���{w/�9g`���ꪷު���\&�ڦ��������~��˹��
�'���W8�O�RE�ei�tI�ı��]��g��ʝ��^e�g)ݫr��+��gq�d��%@�C-����5���n:�|�+W�MC�BSV~hI��+6B��@���%���A��Ky�'�+||��~ϟ�^�ksJd�d{z�D%z{�'O����[�-y/L'Vx��2�P�-�y�}��,Ǵߵ���6�4H5Tb���L�$ne���b�Z$�{3R+I!�z�����'�m��UV������ Ý���u��S3�nʞܬGq��Z5�M܏U�5����%��W|�`�v��<n�����薈k���}_��W�3S��<P6����d�VVi� ���m��.��=����h,�����S��W�B�OP;�`lmCU����뫻W�i���lJM�5�уC�ɿ5�y��gR3|�����+�f�����3\[�?ݳ�=r�}���������']/)���[�fh���Ҩ�M���SO���[��h�W��� ���a%٥lǕKvo�V�P}|������k��n<2�U��S?W��s�����V����'Nd�o> ��(��[g��K�9�L_�2���-H$���S�e��i�J�9nm��F���<��%�W^��\���\z֢z��}�=�IA�{雗��!��
�6����Q�z(7��5Z2\�bR���M����w���X��	�Hާr>��+c�ƭ��L >t��FM�`�E��^�k���_G���J��zs�rd �7��-�Z�Oj�4[�<�yJ�����V�Xu�n��m��ʢ��ql�-"����FW����7�טZ�,�5�,�FƖ���g(��nm�z��=9*}C��<��'�i��mO���di�Bj�q,%т9o	��v��_}�"�JhD}`�_��t0�|S�"[��&� �>�+��W�S歼�C�s��2ç=���q��h�+;!�m�����r�����I6�����X��Ӣ�OE���|`����͂ڝ�RKL3$���O�
��Szn�ޓ!�ם"��[�[S~O��%H�ɋc��'�N
_�M��Y�t�|U~N�]�߉j��;3Gy�;�Rۑ�� [�K�7�6�A�%eu?���h	���^n�:'�5���#�3��+j�4x�F���GG ń��+�5�O8.���������k�o��D2�{�E|g���{wi���,4~����y ��� ��:��/χ L7\�7����J���3|K�D�5ǹ�Ж�gT|�z���x��hZy^�0�Ǚ�u�=��o��~�n@p�͎fhd�j�56�h}�r(���7��}�fRʂ�Ck��e~o�++,}o���vxqP;��U�����ǹgߙ�O,׷����������N�;V%:n����8�asنr׾0���ë�[vd8�����.vd��u�E�K���1y��RH��.�ĩ���*��7<si������wr�I0��ZQ�ڼ���Ϲq���� ��[�4:�}N�[/z/��s�Ӊ�It�dN�*�n/�̻0�f�{O�]ɍ�����
��D��-[6f�F��2��?�>V��'��NX��$�(s�ߥLz�=l�<�6f��#~׾/����zG<|4b�\=�E
]��Ќ���<|�b����Sz������a�ƽ��_9�}����bQ�ѦS7�͟�S�h�;e7I��v��;�O���^J����o�K���͙'�]X��+���?���S.�����H�:�w%��;4J8Q�?y�|���ע�!�&X�Lh�o[!?P�lq�C�Oݏӹ�'�D�}J�9=��</}e���w���}O�};rY�e]�3��l0��Q����}�ޘךϔ�KZkr���Nq2�_z�p,�߲���,�������	'�H��>�]s}��9��[����W��W��On��sU�n&m�������:�g�K.�,VtF{�*01�-Ŝ^C�Z�ރ��5�oH���O�V��t�|�ؒ�woU�>�c��?]J&�=��d��|q�pCV��v������_�z�L�U����l7��&�]�!%ٝ~_�������+�ϾԴ[5�mE5`���뗛��ľo?�m��Ή�į�*?����۱:xF�髯��"����Jc�e���ON�#�������}ږMۙ<n�\:yl#��MΒ�y�?]�,f�1��ʱ͗_��sYS��_1��s�(�۶���fP�N~�4L5��V]�RH,�7,<�����F�&���I��w���AJ�geVӺ:�퇍i½F
�%
Dw$�7��(��c�"M�;�%
��sVT�Z,pqCyKsó�;�N�J�Q�
��J&1�<m�*QN����#�t�~Z������[ڛl��Ժ�R��9���3�c�����LVsg���5�=V���:h|"��zL<I�?X7H�~JpLs�̴\hg>4d�h��3Y����K	��{(a�E���M�6�#��b��	�ܶ��_�����J��H�*�����[2�.�ʝZ�d\�M��,�pƑr,����ˮ�+#�������{��������]|���A@E�5�F�hOE�81qo�b,�.>�k4�G9f��{�ݗC�
��R�:��D��S�i�GJ�56m9�1E�x�tT������7SRJ�x9��hIF����S'f����9T����b|�j�S������ܙ�./�/���O�s?8á��c�N��n͍r?����~����S"@a��]���ゃ��*�^`6���
�S�5\���F�sg�<�l�ݶ�j��
5)s�ۖ�z>��d��n�8��c��@���޸����.�d�"��9�C9��?��fi����J�Y8�{�&�J����9	�iŜ���#�&�<-�8���^����,��Plq�>�lyZ�~�H��Z�-�cm�6+�3�q�z1er��Q�Q�������D���T��kdJ�vf�>X��<�T/T)6\ju	��d*&���L9�;�30��ޮf�MC���mU]Z�!�J��}�-������Z��à�Z'�A�e��n�!1N�)�������� /L�9{�!!�^��3l�Y���.'ǩji��2�ތ��v����X�<�9�:��n����Ie7)�����Ws6H(�f����MY�Vs�¸���a�3�}�G���˴^�t�՚�/w����۟�2�,�qϲޜ�&�����|E��vYtC�n˔�)A��M-�-�5����H���]��`�i)~Gmqt7���;��2y��Ȼ�ߕe�Q�dO�u�p�гTt7����	�B�吗�����К������6*4&
W0u̴j��|籤��(I*u���>Q���+vw�^�u�mlc6�� �M�F)�������em݆��w�#��i�M�F��H��U����e�����FB~	^�����NL���j-�`Z����c���c&���6$��3L�LԪ���h/;LFv��z�}9}���g����$z7�*�פ���
�+��O������7�?�4r@�5e��m��N˦a2���]�?M���1�'�u@J���8Q#x�;[�}~�5�V뇅���WW��R����$u�:yTװ°yOot��^��-hL�<�n��M�Gh*��d��-n�[�Qy�o����>
�b0�ْ+4�B���@q.p�e�g�=����[�lI:����c��;9�i�bI�N;�l���������P�tQ4҃i��$oF��_'��~�uS�}���`&���Mf(��{;���P���gϲ߾��}�t��g�6?\X�L%=%Vkx�e��Ȝb2��r$W�s�G?H�ّ�2��W��'M��i`y����!�o?��3"��?������$��Ӣ"�5�R��]Ф��]-�nl�J=�k��̍�M��d3�:[�4�<�����Б$�7_���������<cf��V܆��P��3���C7Zw5��j�(`�f�d#�N�0{�Շ��֎�*��\��%�J�zu�GD�TFp2�Ns�VG\ԃ��־�c,e�������^�`������6�Qy��u	�_��Qޫ ����{��y�"y��*S�p	Ec��g����7������(�?!�yg�-�����ݯ�����+ct3[H-�Nw�>����^Pʗ��H\"MńgK3zn#<g��$�#��ډ�훇�=��2�6�����!\o��f����*+�����;]/^p�1L���53:���4Ϛ�:MZX�$�D�����	�C5�	�Ő�6�)I�_�A�~��&�~������;Z������I�؃j,#�:D����saN�V:9����ī��J��_�d�|Wj�2�>��mԈ�E]�~5�g��J�ͭ� E���j�ڷ��Bݐ�V�@�|�u�P�nv�k4�:H�)U��G�)�vɐ}��L�M��k�!)8�����st�;Ty����=)�3� �Q/�'V��^���gk��q�B�L����P������|�iG6l��oQZ&�~a����{����w��3Z��;��fw*�i�Kp�Շ�˯��ߋEI_����M��F-�]�v�)�mF*�Z���.�0�T����g��E;�?j���|cMgǴ�ˡ_�5��>E������o��Ye�33�H??���l�i��5�xp �)����?_�F��g*�g��rMp�;�Ln�d�2�MQ��z�&��|��Z8��ģ��ޟ���	;�w����ۆ|`�ܞ�J�d����E�]�_��N��o�������]^�.�O��'h�z��X��u��"�E��\�.r]��U�+Uq���|�xjP�g��G�{~�����O��?�Z���i�����O��?�Z���i�����_rjLL���Y8�q�s{���[g�Pܣ,xGⱑ��wS��iՅ�މ��ֺqqI&{k*=��:��w��S��������T����x�ߒ��~����,��������u����\�.p]��u������U�G�	�#�b��ȓ>~��ӄ�F���1S6	�o�"�����y�>��t?��(&�md��]����2�8,���L4,Mx��Г�ݽ83S��}Bȫ��S�P�|7�͓��V�D�i�H�Ȭ�Z�xTEO��e��,6MU6J����2U�`J��l��ϯ�eU�.p]��,0�?��]6��5��3��RV�%�Wv�;,�\�������̛%�/�g�_�5�1]֤>�g��1�ǉy�B�sU��|��ݨ��v�8���#}�������Y�����br����ݪ|�̌q��k\�.r]��u��"�E��\�.r]��u��"������ �o��gb���Lmm����Jm]�%{������a[��Xm}}����B�b��*�鮮����\	�� .��� .JJ���>~�~�7B�g���.Z�k^����7 i�E�8w�N�g��[{<<<�~~�/�����+./_3�0??��cPa���Ϙ�(� TTT���虐�p��A75����t0��9�����c�߬�����ի��������ׯ���	��(��������S��TWW��:p��0Hx1x0Ix|~��k�g��h��ٟ�;��6 ����64�c�>��~JN�dkk�)�>~M}�%�RU�16߫�||fff�x|���,�4)O/hβ�A�@����`{��A�F�mҮ`�dɻ���X��U����xCMMm�×l��zz.h13m�LG;[��LgG6fZ����[�.�|����Naئ.�677���:WVV����4J;r��\uһ�����V77�y	�_s��(l˶�
4�qiʹ,N�(ަJz������6G+�%�oJDC��i�_�	���6h�52���mc�\�|�zC�J���0�Iǹ78˸^�ձ�E�8�=�N�Ŵ�P�z�ko_�K�Y�~a=q߫����9Ϝ�S���f$l�^$��*���F2���;������LNM]266V6-�wI��XwE ���Ru{;�NU���쯗ҝ1�9��˳�֤�������bѠ��jN��ąߎ�/�"*{3<3���ٕ���Ƒ3{Tda0�1�XVJ-LzI��A��(4K�o%iK~������c��Yk�E�Qk2Zi�%n�p����%i��;���'t�PʹZ�M��W�+Oҳ{�f�:]�;Ǌ�T2�[���������E�|we7ڣ3]����08����}�+�|�����HfOz��8�aw/�ypL�I���;���8�v��0r�`�綱�Wf�~v�|(������ܯ�cs=���C?��O��_}xT{X/V.J,Vh�Q���Mu�~�Myy*��8p�?5�;�F#�+9�����9b0V#����{R���J��A�R����;ev	d�SS����`w�s�����
ܙ�ƽ�lmm����000�6��Ps�I�#��->w9��ʪ�3���B�.IKKM��'��}�9���Z���M���y(�Z�uHPa�����M��1�XĦ}�&�)5�F��^�����lPs�<����N�3u���D�#�@�g�/^����l�cӕ���_/���r���$�R�ӥ��m��$iW�N4���S�u�x��2�\!

���ݢ�q$u�)_��:|����:Щ��S��[�8Um��hU��
�ۼ{�K��D�U�@��/O����XJ-��9x������0�Ϋ���p�̞is�M�/�Y}z�����@~~�i�$�>aR�y�����:E�C�<�B+����-a=y�5�>� >���f̥*x�aa/B�ͷ���vGQ�F� r�h����;�[Y�e�������9@R��?������W�up�r��������E���B�-����Ѐ��{��"�6�܌A��3��%�%��m�l��K�Sc݁�E<����09M�c�8�T'I��{�޹P����~j�����n�t��]O�I)��;�S��F�!ŹRX5���l��v�v{�j���6��h> ����۪h��w���?^WSCe�=u��0��mߩ�.��.Dʫy')+/3������a�f�,((�D��(L/W�cojty�]����׵�/f���$�L��E�~��m׽`Gr��gQ�܌e�ٶ薍ۙ�xf"�>�bͅ2��M�g�n*�,��aQ�U�/�� ��5ި�}/��\/��լ)�<��}%ZN�%JS���{�^-YY��'{����yfݞU"FE=�^%Peq�����~lz}f�UKz��U�I�<bo�J*I֔���i2�S���/w�ªu@Տ���^�����ʤ4���["(��d���0ĩ_�~���ɉ�*�;��<����[�@���U��l7;
_��C��i7d��v�1�֚�TΠM�)T�!�S[�o����H�L�n��lsC����vUH�fnN�Ѓ�O��M�T�����Ӹ�t_��J�����/؛��h��S��~�	KN��ne~��}�>U}�1��u��ϋ�/���ܯ�<�����:��-���E�~��=�2zʗ�Ҟ@���:��J&q͵��܁L%��k������A���wg��g�s��ͮ�Io��.�ğ�*��2�4����e#s���}r����eذ����.�P����GJ�7��I�
�lŷ�$��N�|H�d��@��[�K�DO
���:��{�awF��fy�WY�#2��^�mMK�b�>=h䬔���s.J���fө:E���Ϣ�T}1�3�m���O[��
��i�%�?��D����A)��1��]<��ͷr.������k
�݇��-���ݰY��~]<��(�L����8����Л�n=�[2 �w��st��9JcnaQ1�q��݁)� 0S	SR&X��!6&&�H�k�>}�$����tT�[�y������8�{�bǁ��+��x�F;f��r�U,nd�~��D�N����%D�_�CM�rvn̰0@�l�˫�JZ��Jh����� ��>UZ\jJJѷЋ��e9�Z���g�W�e��/]sS;��h�X!���������xR�COy�PP��|C�H��t�����奅�.���0؍~nL3�+�B����Tc������T ������_s���|M-���2u��v�3�ť�{����_׼�	s-+%v�/��+Y<h��8�c���pQ[�WL0�*�R<_{���tg½���+���v{qU�3U�F��gZ�4`B.O*F��8� S��������������0����{m��������� �3#UR���B��Ϯ| R��A� LT��J	�Ef���^�S�7i!R��2�a֨�▆{�5�ű[i&������3t+o�A%�7gy*��������N#>x��T����S ��Jݠl&ini�g�m�.Q�E�mA���75�:tȴ�`Y�'��;""�F-V�GV�ԁS�kW�������$��eO7ϖ*�xH!)�5�NO	��Τ���(A���3��n4�K3:=��[v@�ޔ���˪}���v5�bl�
�H`�≛q��v-Do���]�[��Ew�!�
r�����ٹ*G��ed]������N���u��ҿ�{�8�HU!$4~����X����%����o������
^�n2����:ؒΕ3�a\PH�F�,+x%.��N!~���*q�hk��X�,���9�KDx�xx�bX�g{�)���O����R@zh7b��v�#�Bc0"�x�|H`��m��I)m�:�A�e��:,��?M���N�x�������w�oލ�9����Y�,�3�M$��Un}x�G_��hG���EE��*-�u�}hT������b@�^J������q.��/Q�8��)���W{�oOň�瑟�A��񘋴X��}�<]Qg�[ס+	l���=>��ZG,���5#��k�E���<-5I��w�\��;s��M�ԇ��vghR⒳��Ei!5*�d}K�YE�.��*v6�WT����wZ�8M��vק��������J�����d����-�=q���~)k�~�m�ɛ���� X�|mꢽV!{��JA�7s�� c����e��vl= ɢ9~��]�N���(m�;�l��2�@>R�#5{Ȱ�vu�QZ@�sWv�%c�|��𸡶lfٖ9��u�MY�Bf+:_���z2ι���.2NŬ��Ӽ�� �M��I(
�D��.Ͽ��tu��Mo�l`�\�d��m�:�%=N�g�}u��+�\*�.�HIkf��Tٌ��7���yN�bQV����1���-������b�W��TLuM�K��_��;�+/�V����VU���J9I\���`fG��ҫ��4�fm��0<R�h��0�N\�BL�lc�H��(T{�]�i[񯒗0�w����|����"M�h��-�&ʹ�X-t:\�J$m��7��!t*C&;�w�}Vܮ�^R��O38��P���D5�'c �A��#������h-�ތ)�]��[xȲ��Gc�����%��<rC"�������ۗc�o��pRU��$�~yJm�'geiD'�~��P���!�6qo�򸼔���egl!�F� ��WIJ���Lt��b3�*����0��r|�u��`f ��`�9 *��w��)��4�R�� '�;
;��Y�"ӻ��R�"WE��g�۲��"`���T,[����K�<���Q��^��y���N���P�R@����=��J;��`�s��~a����{��Q�f��kF�����6\:��[�Nh��>9�����s��JP%��������^�u��寉!22�t���B�Q�M<	U-@<�
���|�e�㭳c]]����$y;&^���ug��� �q���s�A^M��V:ƹ��t������kz�y�v�;�9�^�u~��{,8����B���޾��+<���4@�$��`��.>��� ��Dۇ�� ��J5�~�WV^���*:?����]�\0�{i3؎*�M�Q�ɞ���f�7���X���o�%q�y0vW�SE�NI�>�cjEح\{<��00~�#�E�4�W��N!'[���Z�N$uQe������
�Ri7��^Q���/*�N@�8����Rǵ+��I�B��1��Z����dM�����J��������:��eI��d���,���{R��T��a�1*�%r��3��8z���/h��g���l�%�m��ݹQ��q�0�1�bL]�@#W�L�Vd�i�j��i����P&j��	��({���B!�Xz�=�~�m�U� .�"H��P������`,,1U4'h�}�D���v$�02XS'R��a�\����91'Ǘ͊;"{K��f�H�@u��2wA/�;��z�6	�d���혧`�{]c���I&?��J5ė�E��I>��.���r����΍ahq����Cy�E'̱�xGP̉����>i����!cG[��Uq!rB!0��*戹�*���Ҳʐ�V��رr�*Mj#�I���W1��:�iy�`Rl�UK�by��֐I��fMF�I�r���7�m�թ���Ԣ@�:Ss����:��%��?Q��jɣC6�,�b��)�b��<d6Q�WiA׶�W��[��"c���Rx�Ĺ�?�{R欗��-;�WU�,-���W����@{��t"f�V�7]��Ѿn����2依=��ږ�� w��pKz�VV�M n~�������>V�6[ħͼ*��/lYo�ԡ30�Ŏ-M[}Z�!�'rm���)z/�f�������TȀ ;t͏<����`7,
��e�ܹmܜ�1߭�����<�2x�|;���~U���V,�j�P�����3�$ˤX�c��!4ю�jev��*�����4.��� :u}��*���;.̂�6䦂��/ʞ�6H���>�|皟
$Ȧ/�bn�:ʜ��:��L��2��k�Ɛ`�~�'���O �*{���|+�����h~�Z~���A¸��!�^x�N�}�, pX3�?1�>ɀ|�t/`�vz��s����W���	d��@�"ޡ�]�UYH���[OHR��I��⡂8��THJ���!R �{�.PE����hs�%�t�K�X�y��!�VP�ؗ� U.q��Vu۩�=�
ZP��)~��%�kc5��ܸ�3\��X��G����s8�}�w���Pk&_�%�E�~I���NNN�T���Sa�FaV�)��>�Kj�@���:����H����8A�8��_%0�������˶ ���R���\��?��S����}2igU��	��?��K�uvX�/�y�'j�Ĩ�|��H�;K���+��҈�A�����&���VL��Q|��ҡ���]��o�b�,D:�j���`�T�?���W��rQ����d����mY�_�ì6�S���)���0�0SW��뫫_�ri��5�|�i};r�z*QIO�������v�+֬J���Pq�|U6pv����[�+Y
�0�����P�g"~�#�v�0Þ�fX4m5iO1�`^��[���n�Xd�)�x=#����L���_/��*@`��ǻa�Ϊ���ޞ�a^�:
�f�3��[$l����\�Ji^��,]���dMt��{�˫J��g`��%:�����:��8�@�gF]7"��c��xh�n"W��� ��}�G��^ù+˫��"�Y��p	�J��9�^ ��y������}��$o�
A�3�QYe��A𓸴NW��_u�d�`'_�s����� �
=��ӟ@\������9J�/�*�D�sdϴ�9�P1=?r1�k�rAA�D��׃E����ag(r�#����!�Xܥ�Оc�ը��_�iE�9�ҢJxF��:�vlQ_dp��l�C[�T,)$���F�,����[	GsH>�/�T�R2��%���a�79��A���.&�d\��ᩞ��=O�I��:qC�_!2�F��(�I2�qV�q��zZ������ TW)�e3-G<1+�V�d�ikֿ�n4:�fړ#�8���0Hp2��O����P��6��|.�}�ɜ�zs ��+�#+�#��rK�P(#�c5���%Q}G��F��Rs1���3�h�JZ��,;��̫W����Yє�M{�D�u��ϪE>��\�3]+�щP��+�'Nlt˟q䥅}a�Μ�a7T�]�GJUHuG�X ��Mz�Z�&Z��E��`��m�#���섩�I�K�*�Q􍓮K3��S��o��*�ܤ����I�Q�$X8��uG�y�w,���ϴPi���rR5[Y�Ꜭ���x�TwTd���A> �|ƪ���Ӯ�B�w���?b�d�;P��;Z��
˃�zy�*�X
��]�����`V	���,��皶�9.�a<nu^���}� �� 6Ѝj�qqq�;zy�vxAz"�e<�N#{���2
�H�����Ӱ��P	j�+�<CګM���T(`p	����n_ �a)��|"��VT�ƒ?�\��x��B����� ��Taʫ<dV�	q�f�/2�*�!V%�e��d}�Y/��� *��ɒJ��3�ˋ0#~й}��o5��]à_P�3Bx��1��j�]��=K+;�����X@"��!�J�	���k9��,t��`F�g���W��SIh��m �92�"���������Ǖ%��R��'+U	��m[`}H�*p[Ѣ�*�S�����T�JƄ�A�GT���G�"��^��}��M��]}�y`���@=�Ѕ#��G��"5�ei@�a�A���d�o�BbP�Y����,�	\C�HW�����'�AQgM"O�.�`N���(��\��D �+]~.�~w�_0ѯ|��d�`{��X
����aT�����Ɯ��
f��zG.�)5�oZgzW�3R�Yv����4-�#m����b@��\Ǖ|F�x
���v�=�l�?�H�NÈ>s;):$S��e�D��j�fO��\�D���@m��Y\GG�j6��JBL'AgMەW��emT��*�����t0 �i�����Ge�y/`֍�m��Pe+'�^Ǫa�{h�G��	!`[_6���%Z��@��N/�������-��kpGR��lU��`�n�lx�Z���/��W��*԰d;�μ��3(E"f�a������"Ff,>�E�a�o[�QصZ�.`���gF�	���qz����S��D>�#Яt�ݯ0=���U���j��o�M4Lg��@��☌�շ{5�=+*;�P�����9��o��K@i�Dl�rxNl����~uq~`��ZRM>Zc�L��9�ꅮ�0_�+��ܬ^�N������"��^C+��"��BEn�% �`�n���4X���YM\-!9]T�KF��?Q�D�j�.~#u��A# 䁴�\TrP�����RI�����`��2A.Dd�ΘCyN!*#,,�KKT6�3�w\���]�- gi��5"ՐW�Rk��o%j^!��6���������m�6�>�b�+���3Wj�l�@�۱�뭵?��^?� ,B��h���Q��tb~q3*��ٲ�
\�4&{��h���X)�H�t�JT�-u�h�$�����vt|~���ݹ�AWH91a�>n$��~�@\�����o��X�m"
��DſI+��}��;�aO��^x�`��U@?�I��ۧԚl��W���/7&h�Q��Lvzq�S�{�pZ�l�j9�]�)��zdSwQ��B(�	7R����":����W�*�	/��
��APS=�`)�P�Yl4]�cA�%�T��"���yZ���f���l�\j7�V��'�l��A���>���BZZ�A�0��K��w0SwC*P;��Lf;8��dMO�5DuzJXWx��~2��%1l ��~���=�b�(b��E�N���^�������PӏN�P�]�Θ]&�������#�k׮�r⮓π��c�$.~1���K�.�w�4p�#��O�f�l�Y��$�Q,��ɨ3�f��$�J?	��Ѩed��c8�]�k{{{���v=&�k�Ζ��?����>�p�T��J�/���;׃J��o{��� �Bd��լ�q�v1�Cd���Iim�J�6[�eY�<�Q<��-�b�N�}��s���аi����*&ƧP}����B2L�CI���ݺ�{��D�9! ��τD�����3E��	��fT�k�u����}WX���3RX6�'�H�~2�#������s�:���  KK����]��$.B�&�t`	��?l�8*PP�!D	=C1�S��t��D7���Vn�;)׽��"ĽeZ�<����>�����顐��^>��}��t�&� .mx���p���a�Lm�,iG6�F6j����;*����SJ�����' ���	��tU��o�b��˨'�/�m���k�>z���ն�U�]��Q���+!��f�C,ot<��{螘�G� ^� R;��@�n�yq
�
O�{�8}-��!����1C������fj��U�Ċ+q��-�����C�V�$`|�THxV���G_��h����V:�N)�ݲ��|��x>`�%��љ^�L�ӝ@/�<$ȍ5�҃`� QvȬ���5p�����y �9�VW�K\g��u��8]Xe��j^�o��S��@ǆ͟w�&�ο{����gZ�V34��Ds�6� z�;wrK����P_-��Rq>���p�b�२���R:��XQ�J���m�RQ������F����`Gb]B�����T>S{�Q��h��ÏpZ\0����R����L��O7��x��?}8�#�8�b�����N���C8�����D���c
��j܁���?u"���kѥ��.%<U:�/m$��y������o��?�M��<�ǠP���B��Tx2��蚘#���_d�RY�A=�� ��L���g�3L���}���T(_�t����~�5�����܈UJȈ�N��㶼rt���pSfXt�c��r5F�s��7~��~ ���j�4��Lf?V�##2���E���P�Ox渲ܴ��p��[���Rr?O�E@��S��Vߐ�sC[?BE|f��͖�a�^���_eA��Q��O5�o-]�z@�+IaB�X���.��n��Lo������(E��8��(ۍ��h�'��t�^LQ�e��'N��)q2b��C�ܟ�K���X�;+��디��M���>(�4�+��j�UtDP��6v$Q�l^���b�s�zo`���u��n�tJT�e �p����c��� �Fg���͍X@[�Ȇx�=<�y�l�3��.�^�b�9u2��K3���%��,���yc���ym�%NH|�(�+�ؙOB�,���x��:V6w��:��dc�LW��Hd�c���
Ԕ)�ho�G�IЭ���1�U��##�e�8�|������2lQ籨*�jX�ܦ�X�M��B�� <����{�N�9�Wو!�c�o����AF$�!~9��1�1!���vz3.e�4o���N�6���EPU�3x#�#�����cJ�	�rD�����S��E�$_���d�>���߉�3��k7�(��uэ��D��b�9�4?�*�:���d���! U���'��b̏����`���
�%d,--O�I9�5^�F���v�ޓH( ���o�>T�n�����TYZ����h;�32o�����aM�j���{�S���,�&��3{�p�%��� �l�����O͙�m�j���=�c�t����5�a=�,�Ļ27s$)@߉(����E��ag0.�@�������بc糬;ZX���mo�W%li�D.��s��[�C�Cݱ/�$�;ܳm�l�U����q`J����W��������UR�HC�Q����/�e+�}q<� �W��m�Q~N�U��X����P�9"*;^�Z�c���#��OU��6�ӨC*ܶ�N���¼l�f�2����6�; P��A�PC��`77�����%�@�L�IÖ��@ �z�ԡ�.�xk�M�c�Jm�K}X����CҀ�a�>���7~	��b%�q[��&�m����bv�F��;��vgq�&u�<��+�0�L�J� 9��e��i��o�C䨙�an�I��ڹX�.��:���E��N��,��6:A��'�k	96�9b�:>�ժ��g�8M;wX]B݄8����*gM����3��t|8_axLuR1��JbC~H<�Î[��S�&�=������7�I.��~E�M�O�Kҩ��qQ��C�m�Qi��_���]ѡ�i���#�`l���|�.����V�P"�3�̛�z��^7d� ���$ v�f�m�~�\W�~�e�3��]!�հ�]K#@U�U�>g��N͏�� �o��v�p$"m .��q#�76G���A�g6(_�l_�4�.X�֕��Nv]�JBuC���?�N0�^}+���V��9�ٗ��g�u1��oXO0A��W�s�?U0���(B�u(*%5U���&ԡOܢ����f���:�Z�A��u�C�(2��K��x+,�5�&�>�Z;�|L�X?0��_���U�v!F�X�\H���8.�qj��-�B�B9.�HZ��.tq��S�ڂv�k_���'�?;G[vĬ8d=��ܹ
c ���$w/��O�zN�>�l���y�LP��+BJV��ٶ���Hݎ���d洚��#��6�x��6�m���^����3��!v2��P��EW;�D侳�x[�x���9��)�j/=��h����'4�a4qy�-|��nk��ßSCO�3��1�8#q(Q���{��0�`��D�B�Q�^R�b'u�|md"�*�n��6���A1M@�O |�#AC�Ųݞ䫇�4U��{�_�ӧO��Z4h�Ȩ�ԉ���џ�I�t�ۇ'Z�uʉԞ!�b@���Η�������h$���O+%F�j��M��F�'q�D�F��򀗄��;Z��~���ܬ�: h��w��Ϳ#i:��F��5�F�+�u�j�,��ǌ�q�^<��	Gp��b����:Z�>j��C�S$#���q��>~�Y{���~����-�=��;w`y7څdo^{u����`fF�o��tbJ�Ψs�V?��R��R�Fi����yԞ�A!�)��%���E෡��"k����iw $���
�pd ����w{*	��+�<<w��^Β�Ld2�_�L��e���y�L�v�/�Y]��	˖�R ���hy+�m�J*�3ˎ�N��o��5콳�E��m\��:����K�7
�>V�6("�d� �J_�U)o^�f}��ia�.'�~��(�;w��91Y��ڧ팑c��6��T�-,���~ZV�|�h�9�F��S���D��*u7L�~���o�NI-�iP~I��B���G`�Xs�2���_w�x[CK���X*
?"A�#L��r��%S+�.@���@����+��M�<@aޠ���"�w�(v3�Өٙ�)��}�[.��$޳�3�
�tՀ��s%҉\�QK��T�4���U��d��TJE������X����Xq���:OA�q�A>#��a}'�����n�rN돎�5�7�S�t��K�`�����9yO�ׄsވ�`�)ٴt�q�lQ׮:��b��O4�m
9�������l�U�Aw�р*��t �����N���7`�Z����,�
NyO��u<���`f�۵��~��'d#�ws�w;<'�P�
��8�o����-�d�8��K������޽��������� .�/�ϘtTΆ1�Z���5Ң�,e����젎h ��>������(�p����F���zh��~t�i �"����������p�xU�����ml>DA`2�D0A��C��m�;���0ӯ��^كZ��W%��R����Z��OqOzZ�׿V�|�J\���Z���<�m�#�vK�?�N:8揎0kD�^�A*��!�%Q�?LN���{�1pN��.&� ��Y��j��,[L���B|��+S��Αu�d~y��1r,���z -	xdc��4L���H8�]�Ī(�&���k�m&�E�!K1���ذv�O���|?R�a\�x�l}jξ�;K�Xw�[�{�3툧�D�.?L5���������}���"����c*~j��r|C��E)9v����M�
����q��MmQ���[����!����ne-�������-��SAqea��站��<��ۙы�����P���4d\���_�ol<�y1Z�������b"�%]=�
وnƿ�K����x�Nf�u�~$�,3:���e�9�X:҄�{�J)��yC�z8�ͺ�K�XO�[=�^�������/2�;�:�D�1g��!Y��a�8<�j˿ՔM��Kxy��1m֋Ԋ����-���N%�'��S/�)������@�w�nǹA����sU��6L��6��~ԃ��m�/x��ۣ���@m�N��S���/U�����la,�'F1~5���nA�X����.Q�������{� �KA�U�sd��;�܅��@���xDM�q$�7o�*1��yᾛ�O��`bo��d�`s�I�ܥi�o���[��k{��]F7��,�g+&��?R�+���� ������� �A�X�a�7)&Ǯ,N���a5k�$<�6wu�q�3�3�����Vvz-�z��;�t�>���n�c�0ٴ��c'ԛ?�a�,��(�����G�tT�z�AB�ɸ���%L�'��R���%S���C�%�ǜ1�i�(���������6�����c��p����]@=>�Ÿ冲cE�T�Ie�7t�?(��0LEy���[#j��zN+k�K���[q'�MC(����?��������]�Y��Qx���S�j����<��p�梕9�f�� B� ���K���4.C� ؾ�	�2��{c&T^�{�kyaR(��'$]GW�)�)%Ȋ�C�d�`bY���c�$��}`�R,-��������Zv!?��^D/� ��-�r�ڣ���-��"���q���X|%j�.!H͂lzt��/je�o��400�����:$'GdU]ǯ�B��XS�:Z������"t�h�=��aqv��2�*x���3�Ti%�[��]
�z��UWn^^mfS�-֧��G;,WTT4m��;���S��sP����}D���
|���K�{_�s����X����2m��D��5�]B�)IѦU+c���l�B�U���	-%�G{J��}_�uݟ���u�;��:���<��x>�z��u�o�(v;쫌NH�s����A%0�x���)����t>Rń%0�B����	��������o�uvLo�����v@�����!b�]-�,9�6;����`��d�Js�n��k�u5%�e�3}W=fg��Jص�w*u���N�9�9�軿�x�@��� �k�,絳i�%VV�Y���=Qe#��0ծ�X���J�^�BG�|��ϯ�0�(ɛ]��>=1f�/0�d�V�G�gǕ�N��6Ɓ<V�}���p�,^�f��YM���Xcw�ga�Ի�=::t1Ci�j�y�cRX>:5զ�G����<�Hu���T	'D��8W�|sr$�Ư��bS$y"�P2���V,����f4<fG=�H
��-��m���T(ۄ݂#�����
K:ĚG<=g�'�V��a�6���� �F�s_x�['�wI�}m�8?�2^�+>`
��]�5t0嚖��sp ��_����%�q���j��N}�]O����0@o�h*,�9m^+�aA^��Gs'�� o߀�c�ܛ/\?Fȇ��o>YvZH������?��D��Z�����+ ��ڴ��BERI4�xP�)+�tù�9/���U�K����&�6ݭ3��d`݀E-?�@H�k�"������ةkiF�b�+��"�Q'�랞�=����d�[�(�[��U\�kT�ho?�}��}6�x�Q���?L��@���%aͿIMj}���p�����43.L��C�����>�h�-���RL'�i�����T�MӼ{�z]³E��5�v��2*
��@�)@̒��[X���֏�'y�F8�T��<8��=�)����hp�I��7
��]{n7�N�2�䊠#�`�bՇ|�,�5�k��lf�\���9�ۖ�sc=?��$-e4�H��e{����e6_
vj).��Df;�r:66�fo�lo��QtwEo�>���Gp	ƚ�i<���	�nEc[� ��a���S����7ÒKTE��xv�eَ�Z��
-�w�y���(���Lo�PZ�5�`����ɒ��%�-�#������-���c����J�d�'G������T`T��>o�u��I�Y�/?)cb��B;�VN�n���^��%=.�=�TC�����u�Bc
�w�D�.�������t	*A��PR��(=�;;M3�M��
����iV<x�߻���Y���	+�{,��2�϶���;l��k�.T�*��C/�tf2����8��[��GY�X��<rN�[�V �t�6�d4$xs�.�ݱs�\�85��м��DlĜ-X��ku��Ңb,}р����+�1���/O�����X^�M˗��}������~%U"�����8��!����[b��b�7w�ĐP�h�ƸNw����,sk���ak��s�-w����du1hg	0�$��)&En��W���Y�����]K�VaP��2�YЋ#�UL��<��l�p�O1��[���^�?Tpa�iRqHE���4+{���߇�]ad��]��O�����(0Eg��� �ws��?��H6��Ec�K���J�����p��.����.]��bq��e���w��X���{��b�
��S@Z�.r�o�n��m 8y�/ɍ?C�/ ����l*Bh��u�5�Sv����?/:GE$a���� ���JhT#,��]IQ�;�G���������-'U�`���c��PCׅ���d�'��/AF�
Y�F��\�q�3��v^�ӏ (g�
����^�zjR|{�Ý;=E��:=-~=�6�[6r�X�
�aAᩞ�t�;`K �G��g��*
�������n���ŏ��3��!-H�y.ͭ�\[:&���1�6����w�ӹٜɞbF���[�E��|��>1��g��5�L��Z�0��Gj&�4�P�N@�_Ϳ��?�s	�5�!����|�Zʳ��	G���O��Fv  f���R�^JII�u�V|�,�>,��������ʭ�u�A��LW����A��h)���?�}���ݗ;�N�����"\EY�����2�O��4Â�jT��$̑%_H���Ę+FK�o,����wqq�h�.�5GU��~�|�m��S��/�w���n苙L��~�?�ﵢ_�cX����j�`�#�S!�yE�#��1�>Ăn�h��U�ww����u��π[�r*�"�շ�a�]&�"�����Y������e�������o�
 =����Xה5XR\�h/��
'���: �R~�q����A3�D�L=וX�T
���_u6�N/�r�zޗ�q`� �yay%��)4��yHfN��+��"��n�$�jTѥ��M���4d����D�����2����n�l�6�>]��s� %
W�)-��w&����;g��ՍE�a�H��BP_/_�� )k� �n����������/SB`|�ܩF�R�1bDy�ݿ�鮫�o@�>˴�J�HW7�t�R��g���)���pv���^&IQ�J����̛�0���++W�֞=���T��YEĨ�8�P��٬s&Y�x%;� <��/\�1fk2�h>�ȹ�;S��*�>�:��~n�~nD���c�����*b�5�U�V\G���b�j��|�y�`fn^����J�y��aO��]��D�'�ݦ���(u���)0�
�F{��bf���\���D����R���K [�b��K��h�#��k�5Co��s����������؂�v�-^9̉����	����8���d/&��i��D	��Zc�;:hTvq)�`B���ue�����65�N�-�j���OƉ5)]޻��?���ij�'X4��'��F��a�����;C��w/�Rb���/G���>�ҳ����_1s^y=��9�ȁ�+��d�C8���qFs���h%����_Q����������4�6�<� E�@��K�ZOVc�̏R1����NRY�b^l8�H2f�Q� �fB�v�E0�]����F���G�	41Μ�*��~ z���{$i�y��Ɲ1E0�g�D�x�u
.+�IY@�rd��ځ�����gX��"��%+�Н9�ҍ��rr\i����(��kZ���p2z{��h�=X�$ɀ��[\��D�B�<<F4Y�b��r�P	��1v�6v�kLJ
����_䤝�M%�=P���cYN6��[3맅 SoB�-��8$d��6�����UQ�o��+i�GH�2 
���%2��e5i6�S�����[O�z�IQ��-��������F������Æ���y>$�Yc=��c�;��;d�tH��C��],OvI���~+�.o�`h
uE���4�'á,4���X����S�爋�ѷ�� /�F 0G���3�u��^|y㏠V�Y�Oi��4c�H)k�9^�;��|�͊�`f�- H6�RH��W� ��E�\��M��`|n��K��ɺ�?�I�5��O;�Dq�g��_[+{�P�54�l�}��ŵ5����mѶ�q		~$�*@�wV�!��j�!+�~��Ѱ�|v�6C'܆�����p�2CG��J�4Ao�ƽ-&�kƸ���u�?�)��w� �V�8�;s�n�#����@��M���ٕ�u@����#��i;w�,�&�ob�f�����$!��M�(V���֨)�j�ȥ{r��b�b�vh����ѫ��v�5�*��c�c  TA��L��Uű����"gZ��1^�/����ƣI���%C��<ͮ�ʏ����E���S5����B򅞙z��͇_�!w`��b�#�4y����B��AAAԨ'����9�f^:��@���h���_qS�Z�[�1N�1�AB�Qh���)=��
��W�}�Ġ������F������2胎ֻX!j 	�>�D��ִvW�e;���s�Fr���#p=Iʹ��X���߹w�0��ޗǩ���w���t����L͑UG\̦�����Ȫu�#@ʘ���`�:�
/�jnf&R�����ո�{����v�f9IP�Bө:�4s��]��z8��
,WA �[.|����diV���"�xkt�s�u� ���i�k8���ze�:	]/�(�K]Ĺ!��p�zna�Y<�ӌ�1A ��B���/�o311ѕ��
��ɿ�]8=� �w��c2HH�4�� ��}�A��Z�%,���:s�(�Ȋǭ����f��	�ˬ�]6x�h�����P@�J�h�g�1 �����.��$�HU���߯�����,8�����\V;9�͇�j@Q�0���BT��w���D�.Rq�lj(R��4��������p��{ ����k�����D�
:�96����#���&J2�4ﶶ��7*`��i>9�(�s�)`�&q&�r��+z5n�Z�n���o.�������=�kb��ps�&q8�W�8�����x�(�Bȭ��]�����U"R���;@�|G�ʇm���T���Xh8����U�!�X"�a�'%q�7��G�{�������s3-�C�Nz�����VJ'�����~�,emG���@*!A�ZE۬=F�LXqN:�Y��c!2HOD��c�&k��	������*��e����.>���	M,�G���+�fU��C��M]�j�N�>e��_�͉��0o��n�0ֈ2�ѥ��v�D�w^��؁�`��ڴl��z�SÔ1��.�4SS���ڬ��>�X�GK��@�ڵ��#>2����@�t�X��) > �m^]�����$�L�q� ;^?Sϸ��&�hk��bx���8�v�\�����	=��$ʋ�>�d8����$�R�FRJ.	|�a�:�ũ��:ߓb5��<�o�ϐ��@9���@�T�C�)��v�I�?r��7�9�{�m�sㅅ$��{��z�"�&Y�\E����_����G�N��Z��L�߹�tUq�#Mjj^�2�C�Ejr؜��.��zk��:�eO�MC4(���͟i
@̄bRq�&�.���&X�F���ن�q�xX4��g�#��bf�t���.֑7Z�)�쓔iɃ��Q%���saL� )b�^SPdl��4��U���
Lҏ��;�gW���W;k��]��C��f-5�R�Mox�ڪ*^�lsް��";b���ܢ�B�n�������*^�o@p����k�LP��^%%%R��>j�v`��&hR�CM�qE˹pP��4����2�ۚdj��E~*EjZ&14��Yg3������%oT�kIi-[�y��
�|������ϋ(���))$��E�ԧ��c_t	C?f��9���$Ji�&E/)Q
㻓�O���Xl�{a�ʹ +"I?V@������&�N4�|�O�.�A��@ ���IrR����D�^꤂A*� ���(^��T~X�|#D��:��L��rD�U%�`[)�$�0g�諽<R�a��`��M�������mF=���r;Ek*;�:ͦ9IBԀ$2=$���Ø��ν'�P�X�<}�zIp	��$��0��S7qyψ
�~�
��D� ���}XՈ�G���Z��{a�'��fVV~��НY�����(��e|M�nx�.t;��)X���@6�v���9K�Hp�J�{����J�U�:Ds���(/��̣�	w�o�־3�QThYm����GMR��#���Qdm��;	$�s���_(X�z�X3��dz[0B��Dm7���Q��H��}^��,P��od��"F�{�5C��@$C�(ap�}I� W�vJ�U��&�} �ۜe+c�7��P �H���Z��h\�1s�N��5�f����朱&r��/��*��Q]��JL��/~�>A��̇1 ����@w=;���$����a��:H�gz�P��߇Z���,�*�$+�ڈմ���)6,������D��O��'*v���A��N0�w��׺_� �K�`5�*-ޯ��o��l$כ�.���=��
U".}���}ٲeT�a8TUM}e����̮$�h�`D������;�UЉ��Ō>eZF-tl��G��OG5ͽ����.0>�z�J�#4��T��������1.6�K�Q'���a#O��ы�����tĳJLL����ğ/�K�sz� � ��}��M�v�����vf]��*yg�����1}�t��Km�<�(��A\��F��,-�H2���>}:�]�"���L{�ɾ�?���忘Qn�Ҹ��NH�Y���,�U��t�-����*5�E8��vw�:�?$�`�-+�DQ�B�⊁�!I�\��$�>�n�tޢīV�AT.$}�����??�|y}�`Ѩ NC���)�I%{��m�	�U{{8l K���o� .���b�G|�/vZPU�+&}�		��?��m%]K�9L�~R�b��� ���R�X�O����dT'�}��bi�+7������$��X�^H�Xk�,��H��R�V���M����������L�ъ�0,���^��U`J5����FL��R��Q�a=��N?���N�oO!0��� ����-@pr&}6Q�#vӣ�x`$uv�)k0���� Zؖd��d�H�<���ݔ@��Lğp-J/��B~;aR�q����+���I�oٜl��g�ja����ߔ���Gн�>qi�M}6$�?�;�Zj��1��\Q��k�9 �/I9s��&U�+�coM�fh��^d��Dl�����f��ڍi�g�4�E�4w��F0�����Ԍ_��T���L��8C�M2.˃FB�}�}����gb�ňTa1x����������5w�EH��R����\⴩��~'�Ay��Wz�&�d?Au�����ƴ�xP�x��:��iJ���������X��JJT6�F�fn%��/���؈�t�4�~|,\����ǊL���Γ�P��?��c�Y��5���;bb��s/����?]x9��_�:ijw�X�_�5_�d���>w+x��Hf�5B.!@�ҿ0[�d�
�ӓW�,�+�<�]�p�%(��;�f=)��~ɫ��`��/�Sy�ޯ �aA8�7IM�n	a��0�k�^]a�T�J��#��D@�	n�ձ8�G늆��NR�.#���,q�r\ϭ�s�";O���� ��k&��N�����a�+��,�d��e�Iu�qS�?���ڀ��Ɇ���g���%� �T�`�!�T.�:�n� l�4�-��е�
��OO�t�)�<��ĊV�Bq���F��f݉YDL��痗0s�ki�Ϡ��y9�8�`�6��no��|r����c'ô�n��u�q��2�eZ�H]��k���N���8��Zj�H��Aatd�*��;@���5�V����I^^+���R�{�	�Q�bt���Q	�V��� V����V������ټ������k+���������b�6������a���AT��LUTBBB�c�pq�4���%�J�T?<ʸ�B�+
A���k����$ \��o���:���0Y�?�1[Lv]��cݭ �q���A� �aʝ��0�@RaR��1IA�"��NX߇�0X3;��I׿�0f�5	�ϓ��%�	~���c��T�NY�c/�C���W��N�Ǯ@SW�����)O�h��hc�j)�=��Eʽ����z���6�Kk�T�|||�x�-K��+1</@.!�h:	�JCJU�"��E�f�� �8��m���40Q��7!���1��S�ͯo�cҔ<y���]M��U��Yk[*O.�~����m�M�Ci�&9��$b��xGK�2�B$%%�B�� �r:�(�� �3z_�eJ��yI�|�M�C���������m��L�Qe�6�Y%�i�&p�@�N�LP��V��)�)g��"J(��666�p����^	��YY�nkJ���
}x��%�n��C_�[3�jk�a������134}�?w�	ӝ�Į�n`����`�ПEC�<��gB������x:I�F�)%��Y8_Q�@:i�tŰ�����|.3��9�8��̙��A��NI���C�-�gε����4��r>��y������l,��w41}�7X�4�܄Gp�k����]�[�"�W`tj���!([A�
�(�������!DXwjCp��J;bF
�`�l��8�9����%��XW���^@���\0�!��߮�o�œZ��:����с�o�oT�w���a�A��ra��𾎩ƑA�
�D���9��3mjS�=��ȿ��%�⽚>>~?KP��31�mn�����Q N���4����t�Lue�﫱	92��*1c��/�k-'�}~��_1ƴt��-x���ԛO�?D��&8�O���}�<���wfH]�6x6�I���Ys�y���?�9�e�w��9�Al��
�~�2}ss=}'�%�U8?7{)�A��)�PM�I�,3|e{^�R��*�=�!�vG� d`��^�cv�J��G��5@������88��rAGڗck�z��;%77�ٲV�,^�`t�gA[��;�Fp�`�A7b����&�;U�8��Q%��+�y^"�T|�@ Չ��7/�Boo�I|��G|f�F�i)/>�Z/��FyѢ//�V�Jje��'����\����s�7��n�1�4�h�x�}xo�m�GS��N5���s�(�߼?kWj���_Υ��K��V���������{0;tމ-d�VMM�D����2a_o֦FDl��VR~��a�
��'JH���	_p�����X>�TZ s�.��j�����/@���.~��̋�7(ʌ!�0;�]0��Q�J%�F-�	l�r��O'��GGDDD�����׬�i^F��Y��kD�6���c�J��M�U����-�� �[-�l���~�%�s�a�wL^�C_�u�l=�R�ǡ'U�L��\-%%�uS��]^���گDj��o��/���vy��x�̦����ێ 򳅮�d�LO���?����?�f�Ut����"`A7�ď&��	P�FW�U�PA��FԦDGG_ś@D4���&8-��"3/������Ǥ�~C������VWWk28�w�Ύ�)N�!l���]
!~ڱ��aW��F��	�ˀ�&c4;D�D���r���: ���%�����fj���W=�]�f>���NJ&D�AQ����R��F	��nJ|�:wơ����������1Sz�\|i����Ҥ���ZX��ط������kl���7�䝊4�f��x���m�Dh���t��p4>��tl`һ�­�`���*��g��	����oa[�;b
Fi���;�؁�����}7H�f���=747�9�0ݮ/�x6ô����1�Th��76�X�8�Gs��W�7�F�Op�wE|�o�x'SL�
�Q�Gk����S͂�%l����L׏�H���+;L�XfƝ�����v��3�}��捕?b����w�����=uJ�~A��@���_9H��&��J<A�27�J~���ÞaA����`~�4y�3/`N�`��X5��s�wK�hs�H'���{�K��-[���Q��x��R;t�X95��;
�U2>�֌�H�
#�ќ�1��������ӛO:�wjm<�W�/}���}�zL�jE���@���mX�/õ�]� ��k0����O�'���~�8�!�_s�Q���,��<¢��A7��Iw�����Ԫ[r'�-�ކ(���*��}�� ���Z�:A���+�u��d��J$ɽ
!j�C��f�j���� 4��E�{��{���-�L�I/��DV�)ǒ�YS��z]��̭�����ӯ���ZB_"#�n�AaV�>�}H;��ЧJT�����1�a{>���������7���|Wt;�%�7���2���&ø��%f���Xd��7�`nU�3/�m��`Gg>=��Z8G~{�����8��5&�FQ+!��;�ϙ"��� ���#�bW���r2��Z��}Eh]��paz�#e�7"D�2�/HaR�C��D����xx<i��iџ�B~�HK?2o���/鉝Ɨ\���L�An<A10��0;^�*�DM�����c��z��_�zj���??a��X�j�偣>h&�f��t(����;�
��������c��=���K���?�`Dn���J�z3oTY�sM�qU��7c�����#���x�{<��������~/E��<�y�a��2�ߌ!���덄�ob�>�<��Q�^��<C2��Uy�&'Km6Ⱥ+�{���0������L���;�v=��<�g��������X��i�) ����,�ۆ�}���Bǰ�w=�Q�֫��L�?�1���$#}�\l�����������%�F���-Rъ�JFK�_[�hjy�nJ?mFY�|i^��g��1y+�m>Ǝoզ��LbQ'tT���9�p�|�ҥ�U�zv(HW�L��ȧjA2R'K������C�ŗ���=E�s?�!�L��ʑ,�ڳ:$a� zh2�/��̴����񫊊Jo�=p>�=���Te��s�pz�un=�~<P���&f ���>VF!$�0��Rt=۪|d��Y�vu��N|^����!�d�ôq��K�k������0r�r�U�����ʹ(z(��+����cl�lB��=�C�VHS��l\��n�Up
N�+�
;�V�L���o�	5����"�p��X�4���$�	�tU������8�7��/�����t^�G$����~9�N�'e��o��-5��WTTDm��p��"K"���+�m�8�8.�7�\�U�*B�41a�`�?��1o�<|�Bd���O��U�8l���
a���TЭ�yn���+���g��k_�R���*
���[w��zKuM%��w�pRY��p����ş���3{��b���Q�ZB��X�w�]�g���p.����
ȫ�OS��k)u�o���cN�ܒ������������W"`���= 2$EhBj��~�} �����CRR�H�
��Yqm��`~Z�W�Wo��	C���w_�	�LLZ���`���1����mƃ���'i���Z^�k^b�ׯ��6���OL��?2yȄD��KKz�LA�
�P�7<<m+z~�/cw���p�^|iJ{0n53zeS��UR$1[�7�Y�p�]=�cP�����h$)Ju�L�}�7����L�p�ߴ�=��V9��_۷��ֶ���&���NL���,!i���D��Lw6GG+�p�5H|�8���qG�6�rN��	jf��Joo0�O�>}�Qp ��ŇA�q�z�"P��a|�)�w�������z�H�0�b �7-gWH[� I���]64̰��3��z,g������K!V?�� l|�~�ky��P���٨i�t=a�;�U+���o��n�pd~z�!ز�>|ϵ#����3��&�L���Ejd�zR��TYY��9©u�X�ZVV�`�n{o�ZP�8�鱎�j��*�OE� �l,��p'��D���5@�}��+f6kFrU�띊3͊�-� \�.N�[%����5S�%���QaM#5V~��H��!B)�8�&��C���=Ht~́�WQ�V�፫���mx%�/A/X�@3���^[�g3o����@��PaY�������in�I�	�
j�cυ1��E�]�a�6???I3�Y��'))��5Vo�k&��F?s���"��/?�j2�SWV^�)q��_A���LK}/_�l8nk��U/e�oƨ�.I�|��v
}����UO��=z3�-8 (//U��E�d]�o�m[h��ۺ�W����E�����1!��6�9���.��E*Ʉ���|�i��O���5fziֿ�+
�z�h�u'�>%"�� ��B`4��+�������7�B��#��>�ٷA��B��=~3�|�զ�m4_,!�&��t��Gz8f]�M��׊u�5q���I�?�G�~ML�/f�\�~aYe劺�:�6nw�:��Dp�W�N�(m�\�]�����ש�О�ύ(l�ٝ�ĕ����X��s#�FF"T(z�������U!�� V��oEEH~�R�k�W�Z����N�M�S��f0�l@�wv^���i���ъT՟}����'<�V��Y���a����A��qw�w��L���i�'�|i/����D��(ni���vM�q�`t��%a4T��-_���9�%�K@��V��ǿ�BJ� ��ޓ���z3��@��ں�>#u��{����#�˛]^�|{w��DȞ��}��$>�$��FS�_��*Jݪߕ;7.=��a�acQ�!��e��N��V��J�d���_����E�~{�P6�HĪ�
]�EL�����}�B��$aQ����d�����\�(��}��gO8�`�pҹJssw"�,S�TQ!�׳�s�A�"��>ԇ�ǎ[{���I�+��5�-�K�Q���`g�`ׁ7p*�d�*�sڂPD2�љ���"�3������[�� ����*���ӕe�?��bs�ͧ��6���7�h\�������=���_Ǚ
v��Y�eL0��zV
��鞘U-�ĩ���v ݧ-Ÿ���3�k�㏽9����jD��<���@c��{�_:��Gl䩛��Ӝ���$��0NN�+��!�B���eT�'臏�c_2�O�Q4����Rs�_a�c�E���l�O~,��Ϝ��w⌋�#5�����Ok֮�{'���f��짮U�ߴ���r��l8���Y_�|�,���i>uqA��#�,��X!�f�:J��WPQ@<g��ʨ��Y���~!�!L��ǀ�B[��P6x={���T�6����(;g��6�Ź	�ш)P�Pc��?D}��j	�%#0bg|�wͅ$#���p�(㙄����P�aأ;��,�|�'�<פ*�ƘP��؝��M�qףd@]�/��[��2?5������I	/�:���A"A�H ���`a~
�\���.F�L�<��ŅL���Z�փ$i�&cpmP�U�`ۋ����q{e�*p��6�������ͽ���}[�SӢf��Gd7��T�2"�s��bY��)�w*�������ǻw���qI"����^o�)FP�ŋN_#��V[�!do��$�.���Y�1\����I�����an�����Ltx�|���!߂9ɕ�X��Sya�B0-��`���=�����G�y��%�.&rc�� 5�����SV�"=ommeNK��@j�����h-���֟w!e��Z!�"V]�Bd�m�vV�wuyc>n��a�K~x�ٴ�`� ,��[Lv�D=^�wW'��Y��	�*�ӹA��i� �ga!ݰb�%t���iҴ���foX���>4�"K�_I����c����>��a�t�����hT	�>��_)*��o}}=���@j�-��A���
~�)�����r�T�,e��ѽ��E�'6�!�~o�k�yl�`łL,Ȳsp�(�!�����/������xˇO��#+�Y�h�b���`*z�u����$2�ϔc@��0�˰Ot�Ǐ⨣D�{��F����0�@%uw�~���EI��h������u��={��̿'a:'H�Ѽ0̋[� M ��T94_�8�X?u���pU���o$:���3�X��������ZB?��,�?^�!��U�W{�#�<E)�һ6��AR��������b�4C���z�j�����}q8��`���à4�0��9-�ĵ��x,��H
�nC7�%��Z�<���L�ʆ�.ED��	�Z�ti޳R��LUgN�Ɲ�;���D�:uꯠ]Y#է1��.��1H%?6.������_-�����F�+��ԘFVYE���J٧O���rPA�-���x(0�P`����1��ѱ�P<SL�����
ڶ�� 
����`����Qc�8&������B�ۀ6	j�H���Y�;L�`6�2�;�G�ӱl��L�cӈO��g�����rr���@��J������ѩ�Q2ߛEm���)ժ!�5����@$w�L@\!�q�o����]��򮇿$�L�c-���0��;����wj���Ԭ�d����*!:������Bh�c�����R��̦;��o��ݰ���;���k���RS��?�*U��x�Ԃ��Ʈr
�)�,��1&�����28�ڷ��'�� ��7�R�0|�]�r�����&?�(�t�6{5>�f8:���^*���K[I�5 'O8�|��u�믉�%y���24]�<�(��3�u� ����� ���k1��ly*s�/���G꺈��q��s�����q֧�OY��>e}��������)vU'�_r�xt�u	����;˃�b�X�����mb��w���j�Z���j�Z���j�Z���j�Ok�}���q]5c%*9b�?߇�X-V��b�X-V��b�X-V��b�X-V��b����2�����o3/V��b�~�t؈���y��׺o�x��X-V��b�X-V��b�X-V��b�X-V��b�X-V�rk�C7yL��uڰ���5���8Y-V��b�X-V��b�X-V��
����w� �m��j�Z���j�Z����J<]HЉ/N�E&�m����+�;~�)��j�Z���j�Z���j�Z���j�Z���j��lї������~_½5��Ĺ�������c.Z��׿.����;��)jm������������������b��5�����>~��?|��Y�d��5 k@ր�Y�d��5����kzz���م��5��*�ږ�Kt|��k��<�f?��+ެ���!��.N��]k����94���[}�缸(�ߒ�����������Xqa卤���lO�iK�y�+)Ŕ�Y�+gP�}z���g�{���I:�mZ02�E����u�.��f%ۧ�E�GJ��&KO�5~�a��I����O��Jac�0�۞�O�^F򎰓Om�έ�GW��|v~.s��ۤ0���r��&!8��z��:���-EI����coO��9���c�.r�8E�����e�ů?Q-��x9�����E�F�=��>s��&^"�����cs�������:�\�����l��u���x�H[k��F�f�V/N؋VT�z����1��_���X�7��0/�͉3=חYԴ�2���D��X�����j�������lΪ<X��8r����6_��r戡ai��O��ZTӂ�lmm_�)��w��,�z��tS�y.����̝��q�ec�=OՌ�o��>?�����N|�t�����%��$�a:�t��ٸy��~����>7�_���HW7�k�� M�;ǂg;>�R�Т��7�ו��46����̭8y�^�/�%i�Iod�@~�-�W��E�5nc�M��$o�Rt+�u�l��i�A����jV��:g�K|9V$�m��� R?~l�L�.��/��;�� �o���F�;g6��-�ӧ�'>~�������
�m��)�[��L�2�~�&==]&\�A���'=!>�U���Gt���yڸ�٣�����׀p���Όq��J#:3�;���ڿ}!,�f�y�\'�VK?����t>�a��3�ڕ��W�mH�5��[J��Ţ���O~�ٕ�
[��G�pv
�	�͖z�t���$�ky������b��}ʀ�{��v�G:�6���_��^�{�d��B��7)�m^����f?E����k)�ms<�olf&R�(��I7۫�*��x]m|H����N�뺉6����]/^��Ñ��Φ���،tU�Kv������K�����2��.J�x������	�T�Ġf_�G�^�G�3�}ԙq�������\ⴹE��k��+3kA�]/�P�V��Z����@��>����^J�nW�|���xk�ۄ�YSa7�>}S+9+�E=7#�]��	U?�[��;�u�6��{�+2��c^����;�-řF��11��H��;��J��QHk^���3#ͩ�Hn�=̦�6���nq�|F��p
͵�6C_��9֥ɇW�t��ON���4�O�q��N����}��6����@S�j:v�����+��efw�E�B�#l-�Ͼt	F�i?M�����fI8�kz������4ڞ����NjKuixCo!t�����ʫ�Gw9$�e�?��Q���o�Ro�dKB&��o�O�N�iJ���q��)zy�O�>m�y��ѫ�=,��,}��k���V���A�Ӎ��w�5���� ���କ��=fݍ��sMlF|s�-1��T�6ǒ��.�9��!��_Djɒ%�[����t�4Z�^�8��у**ð��IfJ��;zG'���
>b�O�n}zbRүbbbt{��c�k��-GYK4,����N�h������`[�Ao�#a#777zNK�e�ԇ�6_?��;'Z5�|J�2�1�jp�2F8���Mv8�^ͻZ�k/Gyy���	w���������Gdm,��T|#1���mw��}��;&��{�;̓��T@֯2�%''��p�wg_,
1��IIK{�x#�������Z%SSS��Zm�jj�������V���ݹȴZZZ0�����t̳_$��d��d�}a���Z���=���L+�k��G���?�`r4G�� ��ɑ�k��çj�)���4!�6g����F��2������8{5�󄄄��`���c���읾5�ւ/\�~hܓ����C��D|S���O��*�}��mm>4�T�L�>yy~��V�ϴ���oLA}KS��IB��o��j��WY�h��t��u@'��`�l�!ضQAQqv,ѸP���pL,M4&ԧ_����w�;�LL�>|xmӁ���4��/���6iUf�ո/ق/�L�U��_�:�[Z�,��u��o٧j����S
���1j�qۺ��Y�&��e�5�i� �<i�q���w��i�O��b��;�C�u��I��*�>*y>]k2�u�BBf��_}nx�lYm[[��sק�%��n��O���+�׺�u�#�`�wZ��y$����kv�f��#_36wd���I�ګOO�A��m�l���	ǵ/5��'w�^ �P�J_ۤO���)����͈�^AW�K�b&G?.&�g����C��S���x�Og��K��<���C�}��˫���W�g�ߢ��i��>�笞>}6I�k��t���>�L�������'���t�G�11��\h5>Y���m:��^%�c�jI{��:�[%&�2���c��;�7P�w���i�3�:~��#bbr���{
bm'�sN��q�
l-��ˑ8�86�Sth	�s]�p.�������e��b^F��}�˛��5�<	��Z%[�P�����G�6��}���c��=��r�Z�M�Kݥ@Z����-��
F<I�*�5�'�j���0[	�I��I��0���t+L��=��w���q{�/<�Y�jn��I������P�\��g��ٔ�ՠ�穕kV��r�2{����I�^�,�֞n��F�[��3�E�t5�Z�ͼ���N��/>�{t
�J�)����Ŷ��������I��2��O�4����Z�Lw�I_�*��76f�;�:�a��(�zy[��#T�g��~�v���h,��S�V��{ԇ�N>�7Շf���wG�Z�r��_cl��,CD�#��	�F���5���(\|v0o$�#aw�bq �.��!ɛ���tw�O���m0���E���������ޙ�gާtG���+V��EŖ�rӲ
��ތ����:��=5���d�nS��&]5�V���j�=�9p�[�-�� ��vg�x�4���ڷ�@iK	}�߱x��d/�#�3��ʄ�l���"�C��Go��JKJJ6����4�s�5������XT�����bZ,RŜ��=u���+��G>�~ASfC� Z��ԔU���8�9�~�T`+�Z�B��L����RP�ڕ�J{��N3�e<0bG�ӧ}��̒փ�'���"�B1k��Տ���#����&�<5�q~}z�e�0s^w��������&ؖs)g�;*��3�g��3��M�}];�ӳ)h�䞨N���>ڻ�%,bn�pB�"�Bސ͈�ğ����tv�ff%�)*�g%[�m_�#D�M���i�Spnɽ0/zc1�j8y�XV	O�X|�<RͰ��v0�(s�+��C���5�n������ӛb���%�ҵGN����s��@`��-�0l���ƭ�%R*����g�t�C��D&����m�>�e��צ�2�&6u��W��O��.�4|���qd���>�6�~7��\�S�3����Z�"�����|���ۧJ��hv穔<�1�?o��$�:�ڹ����4
�x���7G��i&��g��ݛtɮϖ=��=E�;���05��@6�K�E���RD�q6۲c� ��Y:���R�w�?���t����8k׭=y���᣷#�������G�f�R�j~���H���HM�R{�ܾ�,}�cǜ��c��}-�iv�q����ܻD���u��n=��uqo�^���)~vN(�b.-w��rI+��Wzߑ���3�x���k
��͢u.��!��^v�ҥK��@����ގ����T��}=�I�#�;'F}j~����?��y7(�m�ל��_k71���/l!���wH�]��լ�<=���	�GT���~���#G�d	)e�nDRb�z��j�H�w?�.�l�I���l?��m�[���I�=Rк�"�F&3�u\Nh ���'`�U�/0ia�����h�mi�#�z=�K7�6h�r�$ׇy��uh {�}�gdZ��^fg|f������L��������Sͭ�v�I���p�Z{����vC@�O�vdXrqH �ؒN
`:���5�96ԉ����2�ҮN��]688(Dּ�{<W~mSW�3׶ Ǐ`�߷MeΦk�EM|��l�ӧ�rH���A�lܴi��yĊT8>3���m-j*�N�4�yl#_Tn0�_KQѺ1����X�#a�h��5)j+��{�Њ����8��B�����QP��{��ro�����0���x�&�N%���,�	mN�8�m77�Y.�a����/7�>���Y�V��^�#�[,�}PpT��6��;�?�U��6��bY3{?b��o�Y�(�����Wi @�q�Y�,��m83p�þ\���^z�;D.e��*��rX{��ޞ�qg�����}��:�~\ץ�w�����-�)�-|uv�[@��\z\��=L&��N�Љ��p�`L�m�1���g�,��mrt��og�8�,G�v�C��ԏ����P�:�d�J���ه��0m+�z}�]E&��@8��-a�������W�tF�k�񖜣�v����g�� * Cq��h�#Ge�^��-��Ϯ!+=��P�U`P�<� P��y��-���v��(V-H&9��xl�Uԉ]]ghf����.h�;w<�`oГ-&��q���I���n�n����壷�{����	.y:M�}�����mHWϞ=7�i���P�Fi%7w�2��7&/î8�h�<�S~9�)���q׮]�N~��=����WWz����b:�~�:~�*t���ם&���2X0M1|��X�x����L�r]�&�Ӣf���˗V-��o�s~���Gh|�nP[���S�� #�U�uNՂ��ګ*F��N�w�0O����s39��,ԙ����\���^�=o��YM�`��d��:��w���#��i ��Ig%�=�+�	L�՘:�@ϔwd�ݧ�����:��E��&}D��':����6�17�-U��)�5ܰ�w��=�Ik��:�+��}����������4��֮mAR�^Г����:+��ڈsv�7�lG5���s8��ҲG�G x������CJ�1�I{�-�;2#^4V�j���B��%�nKV+������~P���W�ק[-�T�Y���wc�}̫+�L�Xԏޞ�����N�r=��{�����{�b��6�Ӌ�a��:0��G���.�B���엫�B�Adk4yӬ�/.d_>1=� ��Zq��/s���O��TVL��	!�pPf�h���]����v��7r���P�tn�ZH8�k����w[�;+�u��-�6+@�uD@!�G�*��[�K�>���T<�#D�q���'�g�߾{��,�\K��ಮ�.��x5�u���ޚS�cgA� 3ܴ�|E���8rğ����>7�����0'���m}zĴY�RG��=!�i2��Q��I��;.��M���z���ɲ.{kRN[Ը?�wf�]$t��:�� �����vefL̄)��~�4�Kwdl;Ƣ����(�s�:��
�6L8��?��q�Omm��sC��,��w�c{�/$ކ_5��ޖ�)5pq(��rF[�b�<�!D�!*��fE��A0+�E�����ή��0+��5���ka~h��bX�������e�`��l��+?do�9(QQ��n�����q�Ӟ��ys�9�6|2!�k[����)s�ɷ��S�n��W���]��OI�yl���M��ʙ����e�v�M����v�����y"�o�)о�J`z�~�+��E�ne�k�Lм�)�v�����b��3?��3��"ϝ�3n޼iL�^/ϦF�[�j��"sh�>���.����wM�\z?:2�����~k��&Єג;�������	���8P�������i�b�6O�^{{�� ��S.����ۧ���N,�?��i��D��4���v��?ƺ�٥sz?0j�-���r�~�����]�~wO��~k��|u�y*���>m�zfkZU_9m}_�z�ӟ\S#���}�L�uS`��C��K����t
�O���+'>8�[}��B����}4�F���^�c09�EN�ܪ|ߖ�{䕹��.u�G���I���{��3�%6�w�Kk9�T���^_���������{:��������^<=|�4]���ze��iͥŮ�5�K��ܖ+����~��݋�A��N�;'��ʾ�ǖoy�k��)qB���S�
~\�H#�_�n���}3�No�������}U�+-qu᪟u���]�����c��9���e��ү���z]I?W^���d�9`�;�H��v��f`�ڟ���J���?�_�SjYn)�(OW?�uN	M PK   �D�X�]B��  �  /   images/e79c4949-80e3-4485-be48-c961657b0025.png�L�PNG

   IHDR   d   2   �5~�   	pHYs  N   N }��   tEXtSoftware www.inkscape.org��<  @IDATx��\	t\e��͝%��L2�L�6]��[��� ���|� 
�>,r(h��w�z�Q|��C�xD���S�"���([[���i�'�>�̖���������$��i���Ozg�w��/��^�Dl`��L� �@.hҞ�]��ib:�cf���µC��i���|��J$��{��H�H���]��`cg��el��SN(S�/��.��s>[��c<�s�^R#��922�G�Fd3F2��\�~>��{<0b1�G��	��L5�	2�µ�u��.�����jV���ʆ�D��pӦX�UW-s�j��F6#�֢��-�FA<���=�:�"A�n
�xm'�n
��do�D/�SQ��B����(S�����z��خŋB���(:��g�Yln7�]���{{�9�,�̒�����L���:�^~Y�*�Ķo���BS���eޭ��:7n�v�r��ɞ��BQ=����l�Gn"1�9o��I�� 2D�SO<�ǟ{�D��\v�c� r- �
V� zz�|�E��6<�4t�ɥ7�� a����w���	,������@AU%��vM�^.^1���@��s�<�:;�=��J��ʐ�|� )NfP�d����*<�$%Q6J��"��P��128��$�6n��h-����Q �D4�v�D�cO�c�ύQ�m���Qe����m$^-����ll�D�+)�611!2��+!Q���^j��H��\T��`P�F7��$�ucD����b���/p�� ŵ	wE�yF1����r�}��Z��X�a'V}ɚu����.1�}����p�k�]\k�C-��p�Rr�>"^�q3v�XFl�Y���6�۴<s)�Q��<@^�>`�s7:�)T���̓�������T!�%փ�mJ�Mǜ9�	~p@�Z��ٿ�k�`�DШ����:Em9f�R��E,C+.��Ѩ	D}�D'v�V�<���TW�faO�w2�T7X_濾���S���r�E��	����o��~�}��گ�z����˨K�bn�Cb���܌�cd-�ռDl�w�t�L��B�EP�/��M����|�>�4hTW
i�[�n�QU�ϧ�H� YԘ�'t��pQ�E�I�Tk�B�I$8��+HS������t�"�0���sp����}�Ⱥ��|���#6d.m�V5������Ňҿ46�r���ڰ��ܳ�*��R)tɥ�b�)��Fn���aNc����2�Ra�����Hӹ���[��Q/�Җ9I�dC�"�qA�v���2QoJ-QZ�;v(�/K57+��5N�����+*�Òd����k��y�6!�Ծ���K��E����Ab,�D�e��w(�h�W;lz�M�`ϊ#���~�]-\��H
�L��^P��G��"�M	$$�4��|�O��M���ՕޔsA��������aeSɗ^���vy^����e�H�X[�"d��>�w<���x�B�T��V���q�ܸ�lT9-�F~�r�'"Q{��G�`.�k)�i	"D���~:v��Oh!�
i:�.N;�|TQG��6��Q�+H)�>gVfCs�$.�̣�0�J�l�↣�W�Hĕ'���A2��O�36&���'1]	B9����*��G���RRV<����EF)E|�N\��8F��0��͛�衇��D(�D��������Kn�����$-Qt�Ώ|ݳj�»�Z�������o%1��<��Z���8�Mg��~��k�t)�ի3Ʋa�f��h��)�Q�;Пco�'Dh'�8��n��F��D�N�����i�$�>N�V3��(-Bi�}�0f�w���|��Ǿ� >�Ɲb��+��
Jv��:�gUq�x'����ehu�%M��F�{�7�R�ƃ�q�5�4��8i,��;t�����۹h�"4|���+�C8���WJ�zD��cH��:�r�1M(��YI��#MC�a���%�VM��ߌ;�H�c���Q���+d|�F\w]ʹ�<��wR�:&�2�X!��䵈�s��ႏ�������tw�aժNl��7�M�33�R��?����q!�����]�;c����;A�î)���
ս@1�"�?���Rl�XNj8��A��=J4]7�Xr�&R�r�E�.��v5V����P���"��$��S@U���5w6�A�T���V����aH�-[���=������?��
z��� P|���/(�ܫ��H��2���2<��s�\��>��>@og�̑�8���X�XbSlISS���cVWcv��8I'M�u�Y�XVT���c_s��\25��J�Z�è���pgf����E�4�bA���xnF{#XU[�$�z�/#a�pl���ԛ���Q
.�<���ex�ŗq��K()�`��غŀO�U��b`W97����Q~�]�Ϯ\�f��!�g"b55�40���r���"�Yb��Ƅ��-g�|�3�RRT��[��n��h�	+����N��|��jy��H]������It�EH�8ͥz!�ϯ,Qc�d�s�qܝ�]h���rr�%�D��&��`��R$w�B���N����f�R)5�U����$p0�園Yp-�Cl�6�ؗ�V�H��G�4��u�������`��kmݏ���$��y!AW�f>R��䦋z�ak�M��"Fh7Bs�(¸H����aC��k͝��}f� |��'�V��sPن���o����b�P�F
�bC����cT9#I�{���Ƭ�"��:���]7T?q��ل�JU�J%��yQ�2�H����gv�SOE%��Ն������s�D}�JI#�}v5�I@��D��ER�q��V*}�K��I����Ýw����c(+�`۶Z���� \>�k5�e���g�jWk7�
�ֶQWN8_j)���F!�Kd�f�2�=����kq|{�����?k�R\�|d��m��-oS�o�R�IIj֠�����G`�8�:��H�ܓ��@i>�$�€ �t��c街���A��'�B����w�a��y��Hb֬E��o:q�����8~:�ЦM��̴�CT��'�X�y���@	�n�RR2z?�1LK�@Ŋ�}�?v+���^ى�ڌ��߯\��t��JĞ�ک"~�A�l[� r�$��� �.1���-�-�Z ��Oз�w$HS}r�O��v�6v3��G���ES	XFo�={KSABx����"̝�V��R����ܙ�n�̀����U�����/�}F�{�֠�� DrG[^��D�VCn��;��l�����=$���c�cs��3��n�۵�>3�����4��'O%�蹩D(.n��I��79� 풲����]
K8�`��13}�̸ƶw��by�2�Cr�.1�"�-���ҥ]^v��;�t���]6$�K�Ȉ�l��W��WixA&��B��}P�1d�1S0M#����a���n�I�7mv����I]�R-\�Z!@�醵g"���W��-Bw�nְ�>�%͞Ƌ�\���
nNG]�(���:9Mݷl����\bt"�{��/���~�e�)I
p=��O�9��9vc��"�߮ۅ/~1 �߇�[��~�#=�q=���F]�8]N�H@U2B�`����O ?��۷DOO �p��&�o~��<�R�
Z�F�*��#)�V@�/	^=<��1:GnZB�}~n�vl(ÉO�3wflC,uR!���o�p�U<x���j,_�_'An��y��2�a��H]��T#�������y��Jm����sϫp��sW��S�� F*��?>������9fD�p�z�e�m�ʢ�}�����h �*�?��pd 2%�ڔf�IY}e��l�1K;1d<��ą� ��={ڈ�P[[�+�����L��#E��p����&����͈c;����;):�͛���"�x�ʚo��?O<�3�s�c7Gk���%�[ݛt|%�r<T2@��L"�;���P;w�Qv��*@u�|9�L�d�C���
r�ơ��T��0��8��=�h��#AJJb�$��~�/m.�{�Ȏ��S�ש��m��̞x�rL����d�XZ��G���q�ɵhiiAS�^�����5��{�3(?�|�
*ROut�$��3���׿�_�j55.<��:�D��E�V.�B����="g��lZAỈ U6���x\�rj���lTmIH.�#�GS���*uof�g�Z~Fpr��?:U��q�1J�|F�E��;��u��f7�*�O
���aÆ��7��q�ۿbF|>����nzR�eR��
M矯�V�o���]��xO�j8�N�L��Ro���J^�&���J�9�J�$�iU����$���3xӥ^���J6!�6T�X��2�<"�=N�����}ɁJ���_ӱ�t��N�D�*����M�V�-G�:����#gv��U����w���تl*��<p v�I[Wה^T�����,�q��\���\�?�<��݂٥J"$�WYZ�7�R%�+�@1�.�2�*�+5�+��H1��Ի�ê,��Pǀ�ڤ"���Ά�]�*�E_8��Fn*e�u���+p�L�s����pԶg�A�޽�f~Ms3�d˵
D�ѓ�z��L0&�'5bw�1t�𰽈"�����G?�y;v�R-S�/jC!�p�pl�)h$�W�����F�U彴�D���R�8�9��Z=�(|�{�?�`�)b4�تƎ�3E�s�����;�YZ��p�)F������[�^�7���7(v+Wb`` �R��Q�8c7��#r'J��͛�16�KьƮ��F"q���i�H	�y���xQ+��u�mT9�RU�z���RffrY��B�pM]!�W��&�z�/R%�D�x�fW*��[ `z�,]:���r�˲��.dph�`��:!2��ȝƁ�Tɱz)���~�R���Nǹ�a���o�Un\>���CrQR�	� ��ΑE|�C�D��/է�
mN�j��R�J�:�2�f3A�rAEY����m�Q,H5#�D��nEh�	�p�Mُ�Ue��TEj��=���?���A%Ie>7Fҙz�H[$>�wO�@:�B���ڇ�s��p�"|�ӭ�����7��sf���B�Z�����6��>�9��Z��_�e��\
]T���$��GJA��L>J�5r;!��(�A�����	&�!�6[��vv�KU}I��l��N��plD��
���<�B��FE�Hp,͞�Q�(�"�K��#P�r*�~�k}C15�H[���$��Sl�0��ǆ�<��ܼ!J�^B\�Iax��ܲ_�f�L{P�r	R�q��D� ���.��R6��}}�F#8B�q�Yg���K�{Y:��3_�z�,Q�i�C!�}�8NIRj^-+C7q��&��'A�&6� s�7���>�Ҧ&xI��Q�t�j�e�n���p�py�������{b�G��ٓ$��r����K�U�KƐ'�:hy\��Cc��P�q�!*%Td��X"Gs��?���熯8
�HB�G^��B�r9b��%(�b4��1�Y�6/^�"����|�T�p?�W�=9-%�r	'���%��O}
��b�>�,���>y2�8�EO�9^��ŕq�!� ���P�ZQE���{Ӝ�zR"r��)B��!��ٓ;
��|���fNҧ�Sr�P)ɕec�y��(->J��PD4�pԎ�=ՃS���*z�mmm���xx!zzۆ�&�����
<)�Ñ�����������׾�F0h�����].�=8NB=��?<vx��Aw�Id�����>�/��h�弖�����D�
��)9A"]l�x[}��r}�N.�E�ޤ;�Jـֆ�b�������6�ޤ��@O��o%$������I���Of�����������'q�ϖ�fFU�L�'Rg�>�{^lڤ���ġC�S�M�EH.9��I$�\U�\�@b�c8<gE˝D��	��ex�i��!~w)��R�uK�f6�>�թ>bS�c+�=�Q'Um�jw�K�T��{�zX��߯eK���n~���dG�n55��7q�c�z̄��B�:���Q?��/��'�w
Q���X�֞mu��$()�R��s|��I#c���13Ǡ�٣�Ct�{�5n�mRb�Pi>Q����ǩ����Љ-�N��H�؉���C�e!ӊ#��M��X6�1ԁj���`��ֶ	��q}�ߘV
�`�D�	u,��q�_A{ub�v�`'s���������)�(��8R�O��Q�OmJ��BK	�*�e'4G��O<�h=�4-}N5 ��d�EBދ��J�U�� [�&�F	"����H�&��W��f�dc�+�*i�E���/9=,�m�ի��B�����2�H�}8��x��Q������0�(�݌���-B��Ъ5k�k譯}�h/C���N���lb/��<3s�7@�������C���u�@�l���o�mR;Q���p?�X��V��Cc�Eͨ�����c�c�cΫ�����c/}��]�W����o{zСe�,5�y�|���|�}�yd(Ʒ۷���n"f���rGy�oشV������Z���"�%ԧ�l�C��5��I�Y�$��ȉ����Z����.uO��-.���RS'f�$vAa��t�1�n��EIT+b���'���?
�8�����k��Ih�ӹ3���E{0���z[�_��=[�R� O�Q�7��H�7�e��+�A�+�(6�=��p#���k�KDK{�Q�t��>�9a�d{=TSe���64` �bg����.k���8B]�㭫Jd8@ʶq`��4۩y8�OP,��q��~��&�VӬ&�Xy�ȼ;�c���<�ʧ�cO�Y����L�=�x��*���Ә��SX��
������[���>TX�`������>[��87����s���e#�޳#O<q�JӼ�q�
����
~ʶI/�����&<?Z�����&�\>��������T������²���ɤW?��~\^Idu����͑��cB�;Y(�y@������s�Iww7���JͳRK�W���5��_C`��L��k\��@����f,�Q?����?�X�J��    IEND�B`�PK   |G�XEm��O �� /   images/f99a6fc2-4a50-4dfe-be0a-52d397e863dc.jpg�w\ݺ6<H� ��4)ҤH�$H/�Gi�A@C�&����t"�"5
қ��P�����s�{�{�~߽�����Cf��*�}��5�֐����sPUuU�� ���4<hNRQS��������9u����3g9���Yy�xy/q]��/,#�YR��E1qIYyEEE>�[�7Te�+ʓQQQ�R�2��2
������G������x��d��d�6�,���d�}�?>d'�)(���О:� #'?AANIIA�	����$n�dԵ��qe�|����Vy3���&���ZV��������e����+ܾQU���704���Z�<���wpt�������}��9*>!1�erʫԬ�ܼ��¢���U�kj�ZZ��;:��{��GF�_������/,.�X^�mm�����������_�C��9կ�����������I���TV��<�O��nŽ-o����d~�6@��'=Ï�դ�Z��kP��Q��֠���4�&'��P6W��Ǧ�"<U�$�="$����|�VS�bE%�6i��QH���Ϗ�v��)���v������W��	�ŪZ(�d&es�����g��@�.��P|`��v�z4T��������t�YU"�~�;P��y%ݒ3lE����9��;Q��oS��1���..^V&X�-��I��3 ?��J&�`��d��c��is�w��D�5����2B�P^C�C��A�Ш<d��g҅ L�J�P���B	Y�$�c�ׯ�:���N�B��r��t� L��o�������`�K�{����
ye�V����zӇ�7�Y��B7.��>��{�淲�;'U1�m�x��G��4:��;�������@X��#�P孄�Q=>�@�Jň�Q�o8r߱��*}ut~�v�8�H���z���(%��êw����&����OC|��-����R�ָ{6;�26��H��K~�S���J&:��#�(��+Od��|'���7du����Gh�j	�i �ڐ���ɡ�A&�[�����dlM��&+x�֢����*����s�J��ӫjLT8��ߟ?�t��p���iYZ���G��*�uǂ��0�e�^a�4���P�G�_��u�T+.}�3��󁡊�c�Uc�'��{���Dŕ��.}7�@U ��c�w|h�l�����O&�}h)�^H��>��4M���J�	�w�c�a��Pهq�����[����&��e3\{��4y�s]�\I0��J��h!������wi�dnV�q	���z���p�����{�Rd����q��D�<�<����'ǘ��<�X���m�e�8�01�ɯ��U��]���6�����ӣ8ǫړ̞4!��1����֙��Ǥ���sW^�w�t�*y�L��	��!��}p"{�v�\�`���ꪸ�H���#"��u�W���"Ӄ����Yc�^�g��j-��R}-0��M0h���(]�iV"�SqCg3���@���~�*�s�k�M�*`p��`��3�;�pM�k�s����L!b$?�>�{wF��
'].��ˇ}S���y���a$�pf��ʑ����!����{�B�"�⻈���o�,w�x��-Z�����R�b����:e��Nі��S6�]ܓ���nks
W	J'�3���.b�6�$P�
�`٭���7OV����v��s���݊��;{�Y������jYw�9`�l��HHg����[T���*�í��-c�+|3˾Yq�e�T�^�n�V��y8	����uu���%Q��-�BH�&�����v����Suk_�ʢ۪�U~T�xB���n;���=P�k�a%4�>
]�2�3�� O�O�&���a�ht��4|L�����!��x���lT��+��쇾�a��'t�\�`���4�c+k�r��}�>*K9\�3*�cN㑱.����K�܇���͘ĺQ�~_%td����oL�������us�7����{�ѓs�O�d^�S{�(9y���8�kW��)<b�gj�㭧S�+���mSGY�U��p)�չp۰���-ט�c���9h���fS�萯yw����'�	�2�MB6ɾ��g0�9�QџKO�ħ��� ��}l��R!����I��)�l��A&΁[։V���ݻ+Ji�3��w&?�	~Bm;��]7����aJ��&����!���{�^�`��XM���ջC��-Mw�	�9�HEЫu�p7�5unyթA84�����K;�Q��P�B�B�ƹ���W?|Dn��?�J��M���1��>��Yb���e���hd���٭ؑ>��sN,$���ÀI���X�璔.�U���/�ҏr�^��|�[�7�g�+����^�%)K����e;�i�z���i�ljtx�}1_y�S~�����~x��|�9�d�}#Bv�p��g�gRMr��nuR�ڼ����C^%��>�Ө�:,��.&�Tx�'���\n@�K��l�}ߖ�k��Ժ�J��é^ ������Lΐwl�3��g,�v�śV�I��η�_6asq{�2A	)�3�I��k>A���KJ��s�uo,��7X�E�7�A�4�D�Suȓm�%��/f�3F����g�D��S��'"�����Tj#pS+i[��Zd�J[���EF1��X���o}#�Cq�����D�٠I\���>T˯~f�HńK;T�=8%1�X�p�K���G�L�a�F��[3*H2`�'z-��'k���tိ�����U��c��O�,�M��V'���]���zXL��(�Q�Vv}C�����^�1�v��9tG�]�m��{����A���E+�{�}pԅ�TÄ+��	[�s������e�@���x��l@mJ�i��R�x~�N��s�RO,ނٟ��w6p�<��o�v	m��y��?}���h*rw��^ ��]ݓ����W�
���G��09G��1��42�@	��Ɵ��(�a֐�S��QOj�K�\�\-���"��lS����l'w9�l�=�ǻߪ�~��X2u����Ī�2���Z�s#����k2��QWm��.�]#U� ��	�G��	���u�/N93G�;G�i(ڏ�9y��_øc�_ͷ+���G�ZJ��6��z"k,b�@�̔^\��|[:�^W�ᛙ�?�1ky`��f��.�N�,ϝ�д�U��~7�zxb���M�qȣ�m�T��h��^w�����8m��7(,�nw�1.���(B��{��L���U0�#(ǟ�ּ������7B�%�[�� �]�Dc��<ne�UfN�u�|�W	S�0X%N����}��|��W�S.�ڪU2}L#�t5�+�ZL��O6��L��.d��t�ye������RZ�!���ގd��k�\OQή�R��{���C��t�2u]���Μ��f�T')h���Lw��po]1'X���gS[
����M��z&{�	M���� i#L�p���h�?�to��	�&�=Yt�%�d܂��[��Am7�[!WEڳ�@�+b����l�.H���Q��\Xjw��g�'�ľ�Y����g�Ô�K�����Tԥ}�xv6{�EY_o\��g�|a��ұqQ��&{�N~�������.'�D"�]�ʣx�f���dѡ�ɨ��(J��j�h�|m5<�Ү�bV��Vɾ
���$����H�*I��V?��U�Vc�mC$ 8�#�i��,C�C\��i!�/g}�R�*���l���~� 7�����[
�s	�W���QW��#O��,�Wl�P�OM�\��0����;:W���5�]�R����"�c3�!���s�wE����2�QO5"�Y�S�
)�r6���'ag�]Ɛ�������_�E�����h^�U%ӏh5�+p�~�qb��yr�4����Ne<e��×��.:�e�n������~z�Q���:��U�&+]'������}��`ΑQ�0q�@�r��V��⫎��'�m�oXP���"��o��NKY�#��[)��ߟ�өP�ޓF�8{��ŽAې��6�]lަ�v?T��#�8�t���/�P>T������u>P�i}�a�݉�2��5ժ�KWL�4�}�PZ��-N����ȭo��)ܧ����t�Wj���=/O���>R�I��۱�?_�w�-WU�ɡvlO�<1W�!6?i��Up�pP|���$wG�ǑvE�c���H�b�
�J�[�=��u5�݂���c��AZ��2[���Qm�9Wm�"z����#{�ua�9l����o�F�F�8��¯�fga�ng���3 �`�DU�W6ޙ�X�a,I3�)��-=���{�L�m#�HX۲��g�a��/O
	f5Mp��"��ˆ�#�j��9����<�?g� _�.�0�Y�a�.�G}�Mto'ss�p<�����*�"p}4�aG	pF�TF�(J?*U;��G�/q,(���p���B�um4����T�D��ZR�*}�2Vm��ik�OY#ҁ��F��>ƙڣ;�w��y^����J$��/�(�2'��>����
m�&�U*��u$�}��DXU�+��x��{��pъӧ�q_;:!����9~K��ɦ��"-�G���h�I�H�	��M�P��Ŧ�����`G��qw`��ɻ4\/b3N<�!�(%g7܌U4�ğ^����[�i��z�u��΢1(�/j�q���/Uvۆ���U&�`b�4an���W67����nFN<N���+��FZ|g�L�n���)>��$�tZh��!��)�7�Y/_�ǚ��`գ��{�\ ��!n̻i�!>�ui\�m�U�T������H����v�U�^e�V�i�[X�J�I��kףs�]�B�?R����z�����볛s|���T)S��A �pDe�t��ٴqt�����'��F�i��t����b�H�&	(/���y}�uR�V�%�H�j*�&u�(��ZU9�4�Dμ1Ͻ%����6g=�6���M=jt^���jc����6z�dK�:3�M�����v^�Y�zPv}n�7������u�b}�BiL��1�KCow�5.�~T��k��s#m��� @�����V�w;h3jH8m�>~m�7�( �A'0q�k/��E�D��D
�0�(u��K�տR��v+k,U��#�8� �Ώ��K��G�H �WN�6�.�����Y��M3W<"�,
GəJ$���l�z`�o{\H@\ˏVT��߲����A:
�~f��ȏqfܛe��A�V����-{C�Y�2!��xe�~&w�%����%Ÿ��a�l�ڦ\��
}�޷��X��JR3j�%�2k��/ e�s1�g����6�������o��Gz,կ><4���=�=˟41��RU^'����ݨ�Nkg:���,]zE0�m�{�3OeM,�}�ѝ��� +��d��P�Q[��^Q��K�旔}w��ATFv]��9y�ܡ~J�Kϭ1ڻF��h5\RZ� ��Np-K���!K.wT�"1�v��ck��`�Y��v#@{hFd�D �Fk�Q�����{�'qZò�*�ŧ�&k(�+�b��(� ��sJ0�bY��d����H�Fȭ���v���b��*x���-�u���p�a�Q̨e�h�oN�� �C�\�|��qL��,�$�#F��װ0�C7dه�YMg������ڠ[�`��q�xL���uP�fcFha25cֿ}�t�'uw;��|��C��"D��z�h���;>��&��2si^����e��_��,έ�xw4l#'�?��nѹ�#�dx����Q����[�	�`���||�&�9���ٻF�$���y��S�@P(n���lAҬ�m�x^r��Iq���*bfb^~�e��+{�2]uxG�i����ᅹ���h���`Srh�X�ۧ��Cu���$��^E����ǋ��Wr�P�GUf���� -#oM�k��)��|�l���څ�����Ж�ٯ_J�ӱ-�;p�6�?M�S�| {G��,��t�̯��=Pq�E��$|٫2�Q���<�2o\z��7=f�cDe�ԯ�c��r��W����SF�p.��y@�Co>p7Ѕ����2R��LY�߾jx��3L�2����(S�k�]H,��6��Ď�AQ��F����(�����oC+1m<�σS^~2P�¨g(,x��
�(�YHp� ^F�[0Y�(u ��)Q�y���`x�a�ϵS��{��IT*T�$85k��K|,)QH�����
U�aMe0'��m	E���1�Kdؗ4嫂�;��#��.���r�T�l _(��>�/�Sv+Q^���S��̊-�B�9L��W����|S�����G����Я����?�M�Xfm����Ow�f�r�����r�P��������+-T��W�9�h7f�up̾��Yc��gl� �?���^`��]�.����d����T_�Yu�HbM�p�)��+'ag��cI ��� jS�_��RG#��f����/�����T������1�y��9W:�g�v{�mq���u!nL�=���<K/�Np��M����%�\�Ͱy��pdʆ�����<�b-�;����$`J�������qgY�	 �-gn�6���\�9Q�,�
QF�$���%�Y��R����0��p9x%����U7�{M�������C�[�r�*��.��O�l��\�h��y�15#�>����N�v���.>��V����3a��\�"��]jʫ�|BQ�\��d���JCz%�`z^���b�Du����� 	���'bm��>��g�Ag���$�9�r�8"�LH�
�!Sn�+�}F��"� �g�7�"�L�����E2�y�Ww�q-���4̮24f�!A�ņ�9�S��z����&�(�yC�� �q:\�F'��� �����9�'����ȩ���������O�-r��S�	 �gZ���f�2��ת�����q��EHXZ�����W��5yF�%��#K����xd�a�+�l��w��;fz�����V���9���֤�EL�i�	<�ζq�����$�-�#��71{�QApҎe��#`���D�%{36,��]�v��|3�%BX5ۥu�W=	@)D�`�,�g�|+#��zMه`.Yr��ӂM�3=�{�񱅿q��ן��Y��?�X�X�VĘ=K
�2�](/�K��Z�p(Ϻ����4�!��ɴz���ao�/�5�C�p��i�Ȑ�����ܻ%��'��=q%jm�S ��p�,v����aC��wL	��[ǧR��EL
�z��!���Ϳk|9fx��#ʶ�u�F9;�;�WjO��}:H�#�q������5��jq�����g��PvhY��3!�����Vx5�d�<�?�3XGI�iojf[�]�>	�x��p$��?��R�mn��� Ф��rZi�e��`�ǦL��'�lvB�U���ݥ�rG���Sϧ�n�������o���}�E��x�G��7���n���և�ho���1��1d�k�g��7|uk���tIk�2�%�����=�V��5�}��.���O�ҠJ##���Zu���j���7y9�,����;V����caxrÝ������+���`^	0S�3.���B�i��f%�Vq��$�;?�r��@hI�j�1l�9��qv�ˊ��]�W����ay�Rӳ+�r�:@h� �A[�:�Z�'xk��F��z�� $8�Q�K��Jm�E���*T��}G2�e��^qkM2$�v�XS�Qz\t:�h�x��E�!�F6 ;byq �d��s/�� A����#a*\�;ˉ������ǎ��/\K�*�n⾅E�`}��D���jZ9��6=M5~TԾ��d������q	o�'FD}����꠶��-d3�!L�і���B��ᙗ�/�M�AoI`=�p��`Cv�X�UZ��/�@v�9���lpڭL�G7�Q,2��&߻)�z�\��������g�f�2�v�E	�|��/
(`Z:K/�\���g��@��`�XK ��0n� �U�*�	�c��I2�����P��,�����O|�iv���:߳sQ���`����P�R��?M����G�t��gM�dyiFS|����(���yqn�M_�������0�L�_�U�ϱ:�^O�O���ɒ�CD洂��:�L��_�Q��˓O�*��a�MC!��13��|9}�㛿e�*0;�*'�6(_;5��2�����%_6�ɖb����o1=� �a��s�₥��:ԏ�_\� ;��	���?���KeU{�����Miu�w�.&��L ��7op9�|��I���C*���D:d׶q�%��t��X�����.�]��4��~��xL���y*\�:ɳ�z�95�˯��~"]��Z��-펅�:>9��ГǻK�=�ijG.�p�d��!�E|~��W���P&�wUfJ$�z��@��)�����
w��Ӄā{�Z�l5��0�;����%���=;oF�U5m�I4=>7�j�����K`�*�-wM��(j�K�S�R��A���UYS;L8;[���MM��a�Ȕ����c��pib`��a��!��Q�p���5�_5U+S�
�:qr���26A���!L����!�!���s&��K����v�;]������7�0Awh���
�:g{��/�V-�?����%1~i�z!�{)ɓJ龑�c�b����
���r���D�֢�k�i�B�d9�L�IWD����Q��8���Q��bUvt^���6A��,���I����|�z�ؾ"�vc0�S������*�`u�Sf$�2\	�ת���������C^ZYhW���'bފ�Oؿ��~�㺋���lTƔjx�<�)�	�������Py5�R+����k|�ح�����T��ViH#�?�5���X�����	./*�F�9����"H�D%O������(ꇢ��A�J��3!F#�v�f�6��6#T�����+��W�$ �`�a�S���j��a����[��YK���g�ϾʏȢ�r	P�	�-5�(���.���mVբe��̓<1���>C�I��W��H�
��0�h����g�F����Z�c��̈)�1�b8P�t��\�K"qH�.���|�u/c��xoL=�V�N��*E�I������X�a������~���#�h5��[s�����]��<��t��gg��mJ~��<���e�u2>�~S����"#E����?���:�wr�EB�։{F�&Mf��#���X��y�]3���ion�"�� U�sB!��>i�P�ަ\�ƲF�R!�n�
�B�����
�X�j�7�6e��BY�W�D	J=��ߑC����Tԃl�R�����gz��T��*A�ɷ���x��h6�S`x#�}�� ԅ�P7���(�\�n��6���}d�7C�����@�!��(�ޟ�|�fz��ç�ˣ~H)���s�w�r�Q�w|���������Ƕ�@k�";Ph�F��C唦�|O����	�q�M�RZq�zN)�����^8}A�)��z`E��!r桏?1��^)ƿ\�㮽TB�s5�>��c���tY��{	��s����9�(<���H>�L,���-�� 52;РK��*<ݡ���;�+���d.�a�C��קB�o���Ӆ8b���z��N�T�W��5��(��0f�V�:���Ꮡ�ɫ�f�>��k� ���������x��kՑ7M�3s2k�Wّ(�@A�kuT]�^���>]�aXF�L��yF���;2��}�6����F����7>�� U(w��j�2/�k��5�GS؋ά"��[��=�BXgU1��Ǟh�pܹ�%��^�32j�קa>T�k�K�����
9PI���Ys`�L	�����F��2b��� �Un��9ZW}�:���m+�1�Q�۷[�z�/�V�������d,!��B�
����L�ml:Ka�N������^�^�E�$�+�������#�ߒ�Q�\(QՐ��kL߄��t��)��/�����נ�`�^�9��r��`�L�r2�V��_�)����*N�J�A����!�`��k@�+�.�����/I<��$�r��_ۙb7����d�RV<�UoU<n,�6{+�z 7,���V����NsA���(^p��<��,�dh��z�b�e��gpO6Y�8�r��u ���J1�@���'_�=�l��V�iWZ��~Ǽ2�k��d��؁/�.!��&��Л�V�)����&�m����]�[�"���Ec
km����>ʬ�m��}Ѡ"��&).�߯�#�o�����]ݬս�Y�׹���=��̌߿��˓s�}���u;|�G�KI����7xӘr���)Q�>C�m	rI�4��@�ݸ�Hd��-�2cQ�Χf�3����%Oֻh��%����iU�\\c��ax&@Y\��&�����^j��h�z�7s=-O�.��)[t�#�f���މ�����+V�s�Vmw֗�C��Uǈ+��|t)�3u�fG�r[�q�V�)��^��Q�z�bU!_{�k�;�����c_DG�2��K�;���i��e"k��3�������8�O�K�v����tF��_`�t%uv��I7u�x�+[�Ꮅ(�0O~[Kr?�$}錿Z=�Q��$���r�F���)����̋��V���	zC����E�6'cșk_T�vE��Ⅸ�(�7e�e1=��
����#�|�B$ �nG�YIw@���{�f�� �$�Lz� ���t�%���é�B�5e
G>s�1M�j/�+��,�M�6{�4'To���6��3�P�G-1�E���u3+��OЗ/+n�R�-�f�4+��v
_���:m��͐?�����M�63%5�����N�,�Kw4|ٯ��1%1o���l�y='�f֣f(�AsV����k�㫾u�4�;PemWӡ�)[X�a)Հ�M�sT�tK�o��$�+�%���#��1�D�`��$>X�3�g���<��>=}N�	V���������<�V ���� f�Z�����CUN\�"���^�i����n_;��׋�J�J� TX�D4Z���A8�س��}���qWc �>��5���b��X9��񼏌�q��G}Kևlύb��&E�	ҭ��n]٠�}H��[-�a��/�![	K	G/���HΣ/��h�t����+E�^�´�7�D�M	�L���Þ���LA.��L<d���j���v�;$�}���2l���q���]~�HXx	)l?O�;y� l�`d�6D<��ɫ�6��cJ\�2'�z���dE���+��?|��R��7/�v۴k�P���P�>z�zZ4�2��{|}�������WK���	��i)���J��V��G;�܉9���qRj�ӛ8�]h	�Q�r`�&��)&GmϨ]�w����=���7m�;�7��R�C�:����e����=z�;wL��7�|܌g�?m�bER>G[�g���[b��<N%�S�������~�o޺�y.����O���@M�=�Ks����{,�����Pi/�o@H��&����y�q�����F�v&T���qr�����EDjaD����8NAPƎ�>�<e +�ҝR�st�wU�G~��)��8��w{�1{����AW�[�&�7�7%��e�����Ў%��	7�0t�G�;AG�'�ěx�ZE�y{Za(��d<�$0\���c.�5>+���l|7~����K����	�5���賡�L�">�`��)N�V���[�'�\�~��^?�b�j��ݞ�32��P~FN�MZ/!z��q¤��g��?uW���!�Zo{�rU��W`�B��:z��Ԝ�❭��ɼ���3�j���"��w��`��\���F��jr�`���_������k�n_���W����Y�i=]�D���lm"�4%Q"[�|��VE)�P���a�,c��YU�z��gF�Y�cl���ڗ&Ṱ2��JE`w��R0�u��Lq��v�w��E���{��;�0���Vs��l�~�|��c�c]M�.���_����;`�dTf�C#��yvI��{���Lv�I�bYqD{mv	E&ס��d,&fO��rI�qxP���*�^3�P�{�f��xN=�*�p����6��T��;2�]���ZI���`W���T'&co�ZL��wdxdO�L�*�	<Û�/qP�_��԰fER�l��Ɋ<;��r�4�ߙ��}~�uu$��??299߶�݄߭��0���.=�*f3��=��%��2�IB����lK6�Jn�[���mՎ��˄K��|.�����%��Wе[��;��c�`�3��;�<�)zY��L�՗�8�no�D�3�ȏ�g��J,~���) �.�.��rpi�^���jam�H��#�2�� L��bڅ��6W�v�H��o}��9<��kC���ק'�	��~���#��>�WU��X���u̦��Nܬ�s�l�[��p�,�bJ{!2��|&�������"i��o�A��4�����c̰)�V�)�>D����f+Wr�Wx����A��2�6�{�.JN8(�wĘ_Jqٛa+��(IǨ��_��E-����?<[�8j���w�	���hS�e�Z:6�kS�<�2�.�?��^Ig)�望"|��C3�ؗ�q�x�6�_�����~��n?��9�u�
�ҧ���5��ƆT��2�X���ݐ}���W�$Pw����b�'yR�tb����0�`�ɿ�@T��=p}���d!� ��ô��!�'��fu Bw�p�	�H�h�}��y�^*����*���V	Ɯ�c�Pʃ���cG�FC�E�k���"W�ط���fʁ���zx��A�������d-�k	6֓�6֫��� ؏�S��Q�[����G�@ѿqt0�����PPIG��M�HxK�~o�o�cX���	�^��@|j��>Z;֍��J�I4�C��2�4Tf<�I���L�07�������Ke�{��$�F��#3۽�Bq�Azq�leQ�t�W�U�I�\���@�ť�C2���H��b�#��ڟ'��-�7�w�+�dS�{Þ����=>3۶c�7l�/��nǜ���AQq��BI�$�ß$����:Q���z\�� ���&9���oW������l�8��}�P�ӭWrs�L D�����֓ܝ��N�vϵ�����s],���F�J��j\<��n jŸ��s��'�#�XJl������p���̀�͔��LtF~>�|������F��J�/�+�]��V���"{���1��&n�~��V������[�?���2���3�lz�2�@��ʕ���X�s��.�7r}l��k�!�dH�����ɫJ�$�R� �!���\�D�`]���Q:��$���n�}g��F�D*&P̟2�K��(����M��<��}��{@���� �f���9G7G�CX���ߠ��S{Q�ZY���t�d\x�k��e�~�\Q|��S$���7s!��K^��O6!��2$�
F��ì��A��w�R�D)�c7��+��j��3���'�2gp3j{�7%�
h��r����W4f|MKI+s<�C�<���|��*�U��W��2ԂFۍ���"��Bs(6�m'M�9a��n�����{����RO�s̪#�PI�R�c�'n������{��[,d��}�C���04�o����\���a�5?ro�`Z0RF]�B�L���+�D�7�#�I,l.�+�$sOd>�bv/��:�+�3d�7Ʉ�]��3�9��=evz�^���*X��s���;-{V$�L��yYҵ��/zi���P/6�J�&��!|��@",�Ҡ�:�3ӯ䨁�/��~2�@��c�ct�?6=k%��h��OEɭ-P�Cl�K�M8�w��0,����*�ɳ3T_�R��7�j���K�ޠ���%�
E#�F��G�-�S:�j�Q�����eGs���= �ŭ�Ӈ��o�꣟
>?^��+*��k�����Q��p���dނ����ޫ:�:/������4r׳�`��>���^}�g��|:<��m��_�}
zҁ^UM�-k9��P������m-Gڟ�⢒~��(���'�f�>����Z^�z����N���w;_}���������WߝU�.�S���A��3��)��5�e�_��+�*(=�����b�`��~�`A���7�O�G���al\Ϳ����E�4+	xa�q���coǈ��Fp�r?�ƒ�Ϳc$d`Fa��[Eki�M�N�{Ze�F�s�"�
��:��Z�8!I+�����T�x���_C��܅�G������H�W2S��F�-H��2�r�}MW�r��2��2�b������������Q�k��Yb�Fe� ��}�oa��>2��wM�)�@o��t����Q0p_G=����.Y��;��}�+���_%�� ,]�a1$��E�i�m�kH��]����t��4�!����������S�9�B�{�rvwԇ�u��P-r�~A��Va���$�@g�h���U�:� �U�yr�_�(_X��( aN��~ղ%�*6���@*�u�����[�-UC��l]@��"��ϰI#K�`�ShO�&�4��{(ߣ,��8�z�<Mφ����$�����Y�܏���-C��X��A)�#%E�e���4
����r̽�*��lJ0�#�n�/�����������S��GB�h�����ް4�!����hUt��k�jR#�kW�@vϦ�G :ֿ���~����o���x(�@��_�E��`��\~Q�N��h���tZ�,��BAõ�Y󖢫�������C���*�m���c�$��2��=�T��v�%�8jWj� %vL����@�/��KXn)���; �����4����o����{�yI7U*�;���Bg� ��G�\+��N��f������5�Zgl�W��9 ��6��XG�eׯ�IKw�*���lU�?g�*A�'h���7��������P�wg�/����p��]�_`lI�tf`����Y���:÷��*'X��t�R75)s�(R-<� ��Z7����S��/_�L�{+��	QW��d~�{�/�����8C�۽�UP�����B�Aݖ�}�|�Ò����0�.��n�g;�C=%���=n��|��\&�V�![J6S�������;t��+�Z�!~�װL<8L=�l�e^����o;:��i/a�_�n�#�e��F�ף�͠K̞�ݼ�����X����S�f�bDl~��%��?yj�?m��?U3��U]��(�v�_@��� �3�`�%���~|�,� ���9K���Å�K��7��29����zI�4a��;P�q�`�ڄ: b����������\��DL8;����>���/�j�M��`��gM��j�;vc��]O�%<E\���Q`����S�"%5��K"ٛ��O�oБ8*�:A�	��ǃh�q�>E4Q��+"xjI@�/rBfI{����t6`�S��V���ʧa%H��d���_4���?��p����b#��I݌� �z���~������+���_�1o�y���m���Z��C|\#s�������J��7��D�e\�u���O�;6���Z.q��!�uj�s:��n��י���JZ�H��ƴ���L0v����ܰX`B:�ro�}����r^r*xCen������Q�#H�UY�i��s���,
P!�}�l7d��Q:�������	��xN�+<�]k���C�N�?J�4t�V���/0������
�G��Fl���q謙G���z�j���md��0����9C���^����OKN�3r�}k�\*w]���A�2�+�57ݽZ�Ff|��"��*����#t��g���	�����G扁eP4�{�U��<���3�[�m�#��������o�����	��o}z<T�����njU�/��=�MA�/����Z�W+xd�d�R���;8oPJ��	^�x@��ZF�K*)��`��c�,`�G�r|_����n�]ė3��e���Wp���t
�}bj�j6��^�$f�/1���Xu�xs����(�mj߭=����|C[O4E�OH�JjЁA�|Rf7s��5F�-�R���Cw������������0Hs��Lqn�0��a8�4
v ���	@*��q�߃�!�y�CI����Ɨ4q�\ft��^1s��WܩQ6��B���t`t >�Z�ܱ;t�^e)
�߅�~?)��BX��j��&gJ�샷�[��NFp�>	x�W�l�2L~ЈzMن}@��R�"�b�� i�nF~iDN��&bRf�3������xS��c2���_�� �وS�����xb���⇬h�ٛ�BH�6��U�7+eTOhXT����� �Y����1n�w��x��=��sP���D��.L�����O���qo	��g�R��_�)����9�	W�4��C��B$Cr�]ϛé��}4���p�i3���g�-Ԏ朋1����#?���6mAȧ��������Q��ܺ��m�C䱛�O.�_3Jb�]��J��P�&�cV�%�X��0�0�֨R�;����l����� :��	�AwJ:�-	�us��?J҇*H�����	��pu�$��Ti���m��y�!�ط1a4Lq�pP�D������?�]�9��-z�ۙ�#��RC*وMz���Y��/g.���Ӭ�^$+����"��>�a�ȁBhzV=ђ0�?/��4�K���d`�8dr�j+a.2S�ǅs΋<AO�9!Jt��86]���S�`\��R�W��G�^=���F??{­K���|wW�Ap��±��������������0ɍa�vS���y�������>�*h����_�F�%zDۿ�M�
b�l���C�{�5�uk�QD, 
D�(�AA������.H��Dz�.����t"Az��)�H�V@�n�~�y<�=��~?ree�d͙9Ǹ�1�9VQQLL�n���p��`窎\�x�=K�A�7.8m��)y�6�W��߿���[t݋��tM�v��ڳS�@W^O��\�EZ6",������ �� �a`ҕ�kŀ���6N����r�8�
�ic���Kqhc.@G4 넾��]jbIR	L">�t�!�o�7W�۔^{�a��GZ�N�m�K��B�2D!�h)����*��4�!HsNE��dUZѿ������77�|�uI'+�k3X��D{Cp[A�[��m>�w�f0 h!I��@�;4!E�z)=��-#-�"%;ao(8�7���j=SD�A.!��@�uP3i\����X9��xyg��	"CV��-�Ƭn���,b�H�1��S�y���l��"�f`����&`�O-�(� y�7�p��w����݈��ZI[�r^���~��� �h8���_��aj��Ͼ}� �&+v�Z���H��IӚ�Y��P�Y���sHEj�y'M����'���@{sF�_C�?|�|����Т:!����\!����.�}���n�.dĎ��_��-�K�ۚ���$\"Qb;M��d2-$}j���o2���Ë_1���4�1e$�bB|��6� K�A��O���K�5l=җ18�22��Bd�Z絾uX�%�Vl�x����޻(&����)�-i�o�� ������kMh�_>�Fɏ�}2:~>*+�Ұ��2q�zL�"����t_����9��D�ͽ�S����ʢ�gr�n��9����5��,����O� Mͪ��
��T=F� �A�@[N��aDc=��Re ��0�$��8Q�n�����`<�RF���i��:��P2�߳��`;	�V#�ACb+���1���c��N�1k���{R��� ����rR����
�G2oF��j*�v�rϏ0���<3�������#܆b?���$x�Q�&�vR	z	�9����4D�_�*������!Kڂ�h��lB�0 ���L��L {Q!=�Q5����kP��[��ɠ
~)�V��żMCU1�h��C-���Uq�l�W͜��{s5���>�V4m�z%��d3j]˓�V>�(P�7�j�̟�,��+�u	9M^�O����c��D���E�A�K���%�i�W ��`i[�/iεo\��[d3pO����@>7��(�Z���p��'a'����lQ�yl����x����.�>�m/8%�Nϡ jߌt��f����뇗��;\ة`��}9���o��șƕ����lOX�>�tv_�_܌xQ�"�2Ac�� )*t�Xv��M�t���CgP���5��0�L�M����8���4S6����S���l�b!���rV~�A�>�����H�����7�T2����b�T�N?~�.j�
~�Z���^�8I���;}���0�.�.]�V>����8iv�M_�����uXC�k�;�Uvzz|X?T
�A�F�7���0�Ƥ�2�~�U���fJ�'V,-���57��]���Լ|4��O�^Ox]�s����Gl0�W�����'�X�z"�c�\{l4DY��=s�
�6͗��W�tw�A�F���fgr�� ޔ�����u���楙Uv�Db�lo�a>[�A�W��a ^�T�~���w��[���X�=`*'	�,Ec2��r��/�$Yn�Fv�6��uM����JX?�0:ok���j_(��2�lv�b+�p��*����#��<� ��{E���Q�o�h�Z�x���0ޠ�}�bԒ�F��XD�� �'Q$,W{ލ� ̎�� �Dl����4H���˓4}�.2��Ǯ/˝Q�H7�[r̦ͨ'\-�R���Ƣ���!�MS����0_�'���UBͤ9�N�ϊ��q������RU�37���k�e�ڴ1q�b���3�@�XJ]g)cE�:}*����2P��)&jv���x����h@��s���s��A�,�䅸�WWf��M�Vs;;b��%��tԋ�whZ��M{�uB3���d��]�` Z�^(
��e'lz'��r�-06;�{�R�-e�J�ۭD���JAX��@�ǮUeٮ��,��,r$W#��ࡧz�f�R��I˯�`8B��<ǩ	�ٚ����z:��E]X1 C*�A���Q���Q��d%���"�~�j)�͇���s<bZgfh�e`YZ��bޱE��l��B&�KI�,��m�˝�~�(�]�3�RƂ��,�fx��7x�=OOU04�<DQ8O�K�m��m�q2�Y�]��+;nv�l9_uԖ���;�U�Q��=v���j���ڻЁƷ篥?�s?�\W�Z�KY٨����6�c��OZ}�Tf)J">�M�7�7NN �B��+�:�ٜ��U~@��� d�R ��$pk�J����X��M�$2�@]��1 U6��k(�R���ʏ���n
,2o�=����D�k$_}��c��DW�b�E�����k��PҰ᥌����-�e�{%{�^����	D�����Y�Rւ�Bމ�Y�1�!0H����7�W�`���V�'�iU�+���E%�]F��(\j������]��R���Lp�pϞT:���*Q�T���ܼ��"Y��D�3��֒���?������~s�2��zBZ�0��4͕<r�m�J�B%B��g�q
�j�5T��b(��M�l��d����~h�%�Bc���}oa�Nw �s��/ �K2�nϻ�[j��VPD��x9��D�����gz]�����������!�`F��� /��9:J��dͱ֥Dqy2��.t���(�30gjG�����] ��q:a�O�1�Ϥu�Ev}l���3�y|E�ޏ4*���EHOX
]fy6�x%V�_��V����6�(6i�X�P7<|sw����U�����}��l���]ybߺ�fm�97��t�>Ǿň������^�� )E (h�돣�0E�m�#�üv2z�3�X�}�� �R��x����Ư�9�����q���쑮���Oz�ɣ	�	S
�r�b��������uxY�CQ��y�#�
����+�C�����	U%��ؼ�VQ�#.){��.�`_L?���ʕ�~Q�"���1�us���NXF���>��Q�Jz�ȥi^)U�o;�X/6��Kٟ��S�6.��
m^Pc�
a<����x���j%y����J�_�~\4"�c$��2�:Ȏ���Ӱs�dC��Ş]{���2��ݥY�o�Vg���Ê��q��*�Zǐ�l:Z�������c�|E8l���E4`z\��`�{���:f��CB������b�gUЉu���o��� ���>�D&%��Ձ=�o�B�����3� ^<��-�����I�-�8d�ez��TOO/�0��&!.�u�����=|�Kl���ټRE�WEW�T�"��e��b��-,Z��~s�KY�G�nTE�یL!?@���L��=��t��=�~#��q��>�ĸ^zn�1����M�o��ē�kt;^J���K�~z��F��˰�r��ɠ0�,O�l����i��G����N2g�̎>%&�n�$����_x�[T��~of��h�ゆ�6q{�D�uO��M��(��;X6�^���J��~��{MU��1v@������X�Z��ު�ҘqKBP˕/� xW�O9~*���OQf�)������p�d����R��S
�R�T~(i͙�WF��@��4��o�MAn^��FB���.=Ӯ�@�kʺ��fa3]����4��e��vޗ
�?�M�������}ac�a6�hߋ�엡>���&�`���_Y�u�[ �0Sޚd�/'�u�,�b�I���L� ��n�n~����r��z5աQ�v`��>���'.5���*A�
CSO��
[��u���9� /=��S��������@5ׇ&��d�k�!K���j U���\�f���Hk�f�>��ۏ<}y�Hze���W3�SQ�[��b�"���E��0ٰ=)�`��W�@ÄH��SZ�Y',Z�
�4�T'lʭ�Kg��]��Wz�f��w��P6�	��M��6˸�����S9��!����?�
�9�Nx�7��K%&��I�c���d��}0`��Z���rx qm�Z�"�38X���U�w��ta�`�}SH�û�.��m��_��q��5�d}��������K S�xy�DJ�3�w�AhΔl�8$�==�<s���ڊH3�[n�a�O{3� �� ��&���=�r��o���L��tY�|���m�𒺊�nN)L2�B��7n"L�IfE=b'�o;�Aq_$� C��q�z��&vC� W�����g��L�5.Y�O��K�,�j(xU��o(�v#Ϸr����]Ƞ3W�ש��iowc��z3��J%~)�c6NA�4P��֛�Z"kM�����J�u�J0�y�ud�X�� �kc\LY3��ss�)p�р��@�w��(7jo�h�����9m���÷n�6{�P an`>	�r�ڛ�U%���#�T�?3*Mp���zx5B'��K	@3��]=���_�"[C�D��0��ZL�B6�0Mz�~���������YȒ��� R6����+!]],�o�h;��9^�S8�}R�&��?`��C#�Dx	͏���ư�$�(B��u������z��g�.m=�Ҩ��T����ƙ�2ȫ��$�>��xE��"M#��b^����eo2�p����p�0�x:6�S��1���=�k����ňG�U�P�F��l�qЗ\L��z���zk�t��uE�t�l�)e��$�ÞH�a�N*C/�	���l�[>ED6�}�ڵl�?�hu;[�����F�D���1�-������
lq�^"<RpБ�x���2z�Ma$��X�P$w�!ߣ'�V��b����g��	�巘�xY�nU�e��E��ޤ�ݏ���%`�����-��ݮxУK�G�\9�q\�+�ܽ�}I�0�n�_4�Ǉ��"6�9Y4�����Q�C�ԫ{������_$��ī�0�c�,������9�p�)��W�y�O��V�񄆈]*�8����cA̱�]�oE�y������vɴ�]�4f�?�j��[}1�����)g��#uى�-;��)C��s;B��1|�YTC!�����?b���{�}���_r����{� Ც���'()O����eB�NAH�܈u�c}�Gܔ4z�'�p٣��%,���)���pX�'�ܑ͇be��Z�0E����z�	B�c�ى@�|���G�@�ls��*��=�*|��K�t���Gm�=:�g���Α�~E��59����p7�ϖ�=��3[�Y��ou�V^�6�/�.=�~��3)� [�>��O�a��Z~���N�t���� �s"�0;k�N����Z����@ I���x[S��m�B�RP^F�邅	�yǈ�� qK����#���e�u��Cgn�h=5�y���70��F�4w"��H2H�ė��g��� ��G�7���"Ȩ�]̜	eOOܭ>O��I2{�R����(���&U� �!p���=d�M!l��ώ�L��f`�
�D�Hu#��G�m;�~�^o�08ٮ�p�{It����:�:Z��6�a�>v4G��U���ᡫ:u�vV�lY��;E��I:���	��'���_��~���8 +��2���-# �u~
l*"�{�7� 4	�**��X�j��2�+2?aϡ�,��5z��YOO�F��gЋ�J0�S�is�8|EZ�r$�ĐA������`��W;��#?"ܢ׎�H�b�8��A��D�a4i�:�����M{�"���K��7d�蟢���
�*�Vu�^�|�����s��$�������*�m��R�\���4n�ԗG2�
{F���g���Q�"��O��&HǱj�ۥ����+,-W���+�Qc ��M����2h�r�r�_�K�i�} d�CL�9�&z>�D��;m��/K���E�y��\��E���vL�)+�X����i��Y�������U�RL�g�s�
FyCջܗ�:�Il����ɔ�m��h�U�����$M���f+�2i�~ҫgկ�ʣ
�+z��a��o�-��$��.ֳ���h�Q�o�L�s�
�ms������\5\D����ABNs��3]�J�9�m{�ٮ��v]�;;5
�=��_ë�t{ ��z��-z�C.���p�7թ���1��:���8mHY������K1\Mӣ�'���gz3؇ZK�
B&z��?~#qY�2����޸\�Ixk\5��)�;v{��Y��
�d��X�c��̓�AE#��l�f��a�,�Z-8��.� 5����q����e���~����S+f�b�k������Y8y�VtX��Ԧ��:�c� @c��U�8X��`��{�����At�5�Q���$���&E���&,��x^3~�����;�t���[�5E���KN�K�%���F�(�"l�E0q�:��R� ���H�	�
��=/^Ci�0G!��&�[��f��w�~�~���)r �~��u`��L5KB���gFm9�'���ɠ���@c��9n������n!��fe��q�.��'�I-��G+�٥�����*�M2�4�ב�b��"&��_4>����ސ�mŇ;��8�P�i�#)R�]��ϫ�5טb���$��j��.Q獏�ߩ��P;�J�����V�$ʯN��w�7a����) \2�=�K�)�����7{m=8�����=�D����o�>�ב{X���v��ZD}O���w�Rbc�G�s�_��JnƆ�[������t�c{o\�} _�.Q�M�".0�~��6�7 ؞ћ��r^#�n�׳�s��Ic��ۯ�2{�*��;���-;�����*٘S"�
���
K��T���K˂�� 9���I��ڝ�e�5�T�,&�[̐�ߺ�_���J��d��.|��:�|��뻑�/c�ei�دA���tf�]�b��޾<L]��x���O�zܟ*M4 �W��|Cs�o�����a-�3c����=�+.&��~[q�A�9��?"L�#U�������),[O	�ł�����>�j������mBO CC�+�����AO zf�@O�|�.�vR�PY6��C$�݂�8?V�{��b�O��ڪ��t**��}��L�p���n��{�U�I�Y�'�Nˇ��G�c15��K� �M��\�89���*�A�U`�	�X_E'��1Lsb|��BmN�7}��[�K� ����F�����Z���p�"�싉�T���,� M-[!�d��_��8��6��^efm�e�!��A��ͱ�T��ʪꇛ�4Թ�=O+9��*���-�uBn���:'����7�m��E7�ǯ��+��0���)HB����Uڛ�1�T�շX�Md��-�)�خ̋�飳u�$)�²��a��>*)���x�C��JU�v��6F{Dx]3F<R�����9���Aw*��b�
f�^�놗D�fIJYJ#������:�aK����+O���KAk��V��nI*ܵ�ԵFÃ'�����`;�S��#v�J_�ҁ�<cu�Lx"7iZ !�|��$D(��]u!�7��W�DY?%�b���i*0��7�,������=o`�.̓*}INf杔�A&�H����U&O�ҫ�5��No�O ps�&`� Z�҇�[��/����=<��pn�_�*�ؖG1�#z:�.�L�7I"�F`Bu�v+�ٻi��N��C5�����N����	1�`2�q�8����[�y�-�u7�	u�y�/�C�A�L �w_��ٗUF% ���:�;e���ձ/�P����I��[�h�Y�Y�����h����dSq�����C����8^��C:�疒.�>���DJ��9B��Xn���s���VߪrZܑ>Wֹ�J��@�]r�;�1=A�qf�\�~�F�2_||"&V��(��&��q�E�&#r�R �J4��0�'���=���o�ٮư:w�fP�,� _��36�8��!w���Mo�l�j��H�>�����t��y�&�k���0���Q}�/�Bt��:�d�R�,	����gpOPb&�_l��1��}�	M}F#|���� k!dPWh��hK�Aj�!#�q��h{�CR˷I*�'a,�	�N%�n]AM<}�~�@ܒ�s#�c���*}�k�Z���Aa�Y�Y5>�ă�`G�����?�^-WKE�*��*^W=�V�d�9GD�.�:��ມc������,��&_w�˧�[Y�m%��}U!��:�j(�[}`��U��H�y��8x�V�mR��nNV_hm�;aGk��g�y������V6�]�U�9-��նf���i�"���m�����"WT%)!M�%�||��ׁ�K��~��E$���6���קw���|�@;%[�����4bց���h����I�J���\��Mψ7��h�H��Sl����5Ulo�.L�Y�^
Y-��� �=fS�M��lu���?-Ct���'v_V)�k��̥�FWs?|��x�5�k��7�d�u1��i��U멪��Q���M�?�3��3�-�)*T#�S�be��-����+��p�/���e3��s�P�	��k-i���D�o�u�hf{̀z�IEY%�6�2�`4��x��P�p]�
_��9vR�nظ�U�h�	�_��6?���H�?R��8��1a^��A��T���A���~�PJ\���&���8�D�o��C>ba�z�ؙx�t4s�n�����+;��7<w	����gw�]��K���j��?��ڰ�dCP;��ӡ��k@k�*&r����>�((��B����oR_*)?��gc<���{�j\��B����v%*�lg�[���JuJ����z�/
]O\0I�1���4�� �\�n����2s�4fb�0�N�3���7IV���% O��N��A~�껑���j���|�y��4��LW���LW���� �e����L�*�E�I��MpQ��P�C;P� N�%:x*�דAN0<=�&gf=��h(:\~q��_�u���^��7�'���#q�9-�J���i�9 4�<[7[��|�k�����R���ܔ������-#��f�.��r��P�+����cc�|�f�5�ͩo���;�߷5�EԜ	�a��:�/aʯ��=�yI�V��}�����Ԕ��p��AD��8qF�����1{����,^T��F��I�V����V�/�o��/h ��-)̔>>��V�G��c�?�N�;y�<+-w@�e�w�5~AYU �4x��A�]��B�25�Gp�GT�����Jp���{���}G�y�{�#?ܞh�!��O c��uyA�+(ד�o��lV<Z��J�(yC�v*
�z��}��ױ8盾a�nb���Bc/̙C�"p�wx�,�}��J�j��O���9�*۠�S_�jN�_H�sR%P�x'�xO���#=�i+f	��)G��2���֘��j��"��څo��L1����~	59dЭ6717f�Z���	Ǘ�|�>�[y} ���%���FI�l�I���J�w�N	\���Jm8��,�k= �ZD����9ii��m2���xp]���N����LP��J���*5�:킧IP���b���Ik����k�",��sW�ֱ��:��(��7W����7��Wp�Y���_�A���c��]�v)m���e^�ABn1oEn&�D�����}y1r��♫b_(O���M+sk�D�Y2�3��L�o�@�����>{y������;�2p�zw�2d�A�x����n�g���EGZ�<3NJ�����Ƞ:Y�J���"W|�o��k{-���\��Ӷ�\Z��_s����̼[���(+Z������_)YY���;P�F\�*5r
�TF�	�=t^Z����˲`�)��S'�EgD֞Ek׋�m�����ArcG�>"��[�t� /��V�pm�����S�U���P�}���J���c2�Nǚ4k��`$O���b�0����R2ɦ�4h�̶�K����[q��3��(`�� �<�'�P�÷74I�-���~�Rʳ�d_7����3���'-�b����Ns�����ޥN����^�M9�V||�'EҒ�VFI��p�n�H��-�t�R2��HכHq��t)�~mvH��ȱн�����%����븥������gO�;}��jN�;�_t��5G#��`���@a�کN��.�}4�a�$���'�����Z���o�y*�WNm�9[�{���I�^�5��U�vG1B�d�4ά�A���u5xR��@�\J���0��,Ϝ���.�Q�}��\*��E�4r쉸��/��f��dt,l�1�݇�P��!�?����?e��2���Y�y7g0\cMz���<[-ʗ}��gVo��v���pMڻ�`p�����\+�b*���u����u`.ss�S��tҝ��[c�.L�A��Z�ܵ��Q����,j�<�
׭�F+܆ѫ�Qɵ=�wcz�7X,x��'���n��5"�d9��@_�`Fe� S�(�g3�ہɻ�-*!2(�Ȗ70�zT����Cn?�[��+&|�K=�˷zxfQ�j�[�a ����U���~��r�{CY��suS����ߜ��, !�=�)~�1�n�rg�;��8��]�3�i`�o.��Q��p�5����h҆�*[k����CdPA���c�]؄�J>)KA+�̞ź��ɠ��/�Fw7�13t�=,y�f��T�$}D_ZP@��B��V���YY�f�`�l�#�k���x�V-܍��������]C��.�δ$��v�?tob]��"��D��I��f�nP����:����(��o���2#�EeRʫ��]��K2�.p�6�L�A�tW�)����w��w>�Zѡ��ҟ_j�� �	�!�k��Y���� f+�%Em4��C\edꢓE�X}܋����]|f����b���=��T������ۚȸҐׯ�h*�إ";߭����_{����N&��������ܟ��>��O��U��A�P2�����O�NQ2;�õ�/{�N�*��ۢY|pr�|���otT'��x�e]vJ��p]%��XC�L�Gc���3l6�ߝ��j����Q�V����ʸ��{a�u�#u�ɹɻU��J���nάa�@E+~i��*x�ܖ́Fg떃���߹�x�/�)E�E������> �)$����d��d-�v.FH�A5�]]�N��!	�DE�|t�����z�@�Df5]�d���Ի@�$�%����곃�c��ʮ,ˏK[e�]D��GM"85�^d���4��y�����%Q����� �fcy�D�MS<5�j�����+��LZL����DQʬ�gf~���x�`�4���� �g4��p���6�<
�6V�gg ���*�ƈ�>}�$�2#�!9Oܱ="�C'k�:A�)����E�%���u��n��A���D���6��ظ�A���ʈ�yaY��iy�j��7X/^���\�y�`�|K���i��<�:o�dl5�L}�Pw��<u2��h��a�*����Ɇ�7
DU���V�)ʠ�Xb3*��i�	;�|;��E�����3���1��K�I(�c���&`��ɠ�=��-0��So��P��'���>:��?�`��^ڞO���N�{����	��"�����`�r���/1��g��AC���O�A��8c8[���G���	 PcK�v"�$E	���G���_-0�:n`1��j5Gd��G`n�����2Ӛo�\6Q�b�~J҉�`�ÑA24�����E��S5e�Z�'ӹMQU��ׂ6#�C�\8�7��4o��-*�0Z��r�^�u9)��6p��|:�:�l]M�;8T�.f��/[����m��z�������������{�<M�˘J_��γ��K-���Cm��1�*D)��iwfR�K��"����lz�Q�T��L�oDW�o�O����i8ƐբL�vUc&��.�cL*՞�h=ϓ&���j�}����̕75�K��?����g ���Q���M��4Kk�I%��Y-�(���I��d*� �K��X����PK.D����CGW�Pm��yy�k��)�s+oW=��6�ZI(��>OxӦY]������g�<Ͷ�]U������0��GX.�_�2̈́
���7J�5�k���9�ʃ$9\��b6�1�7*�
��P��#�D�OI�2��kD�3� 6FD	���C�A���ݕ�0�nR�@�=��&�Fj)p0 o��Fߔ�f��<�pP�;��U���x��AV$\>��=�-�	K��y�>�i�ƛ��Q3o���e�k��'̒A�����J{��$��;>��(�t��gB`�9��Q�x���t�;�O:��l$Vn2���K�"O@6��fr"ԷB� �h;3�g����ǿΪ?sV���c��wW+ź���M��/^���G�X����hA�ba{���Dj|l��]����#X�l�.v����
��o*k���+�b���\�[Y�T��Ѱ��Tl���	ݜ�n>�9s�"�n���O�|�v �p޸����c?�N����ق��]XjqSuY��Ge���Z��'7�N�b}T}^1�f@�dZ�*���	s�w����/4P��~�J�h�-"rf|iSZ�๚�_��I�^��8��r#N((�����SP%C�(#%�7�$�	����T�Yс��VNi�$1>4�����w�yyJ]�2f��ٞ�՟��*�`�-Va���;��U��?�M��0IQ���2���a����P~���eO��һ�J/��7�=���ӬQ9�,�V 9�$�ӟ��7:Ak�$ �+F���v+��� w����ܕvq���]�$�޿�����>D�Kg6��L���sܜQ��g8�}�Im���Y��2)uW8,�,W��*��QM	0��哺t{����8������B���͸�d�3�;�).t% ���J�6�i�4��6,���V��7V�q0�[=?�Q��U�+����2�b�� ���o����Ay��>���?bwP�ăp�B<ȠGdд���B�+�"�R��5�5oJիwk�{ɠѻ��� �$b���Q�z�-у��R\�~h��!���]T�
s`i��Np#�<sH<a5H���ֈ%�$b�1��f�{�R�a���"F+%���*o���	�(G��p>�t�]Ɍ�a�xK%�����A}�$Y9�)�g�Zl��u�'=)c��1��=	�Ŗ�?��R}?��Ra��x�z�eR:O�J�lQ=Xϩ���S>\��7j�$�p��F[*�2��Q�G�
�3.�Gh�D9ǫT���yx��@��oh�	0����u��g#�.(Ѣ�0*�"Г�t�`�c���G��������nRy|$�/�|K�����K�j���tj��ȕ����l��.�?4��p�s'���3�ſ�z���(�>�"�4�<8�%x�}��`�A�!up]�D��}I�Í`�aV��[��^�:�V��.>p9�tK@L�C�S��Gu��s������;h�V+��g�^�s���k C�8���l"�c�B��@F�1CaU�3���s�,�qr4����.�\�%R��A��߽�}���ը��:$�B�麤��І���r�{��m=03ϰ5B�9�d?�t����?{��5|�xO��҇Й���8��;eI��&�ZRi��/�}6�t�B*e!��	��A�Kټ)���ЍwL,�ۉلG�; �W�SaDe�-�t�Q����{�"�6�%ڬ����R�_�u�D�})��BS��f����cা�{��qd�ͻ�����Vk2�[�-$�<�������K�,"���?�98��z�W��IO��h㞢���}���]���<���YT�Ĥ���q�0].�G� |]�juD��~aj�D�,��4���*�Jj�|��m�,ҜU��@	�aH6���M��ƅ�L�pɳ/��n{3�9}wYp�&��2��w��3�
(���ݣ�lJ�W��(�^(}�����S})�|7��.�$�AQ���s���%��7o�5��?3�O��=�t�����Y�b��1��m�xjCNq�,r�턚)v�%����u^�u���@Ǌ�mYq����>׾#��5	�]s���9O���\���q����W1O��{f�Q��e}qg���hQz��h���|�d\p��-v�};2hy�X�/�"���¾�A�^���b�Q�Rz��*�8xJ<m�S�8:���]�奁*A���Hi@�D�q����n�*�m��:�D~\!�T���S���7i�8U�#_i�{|�K�r�Ҹ#C"4�����tW]|��I�3ꪢ&M��I�I����e		J�03���;���&	m��iV���7�Y�G������Ȥǟ��!u�Z��h{A=eZ5�Uy0v!�,MB�3?�TWh�^5!�zjf�	��r<�׀ڎè�#���K9���L���s��h�9L���ѹ៓t̯��<ҥ�>���U��6dR�au-"�!�iL��� U]�w�4>�M7�<�Xɝ�~}e�VC�~��C�t�䎗���B� ?Q����ߔw�_"<�����RK��j�(i��"b��j�i��%I�s;�&F��)m��I�Jˡ�n���p1�,�rm�fxwjvƂT��&��w5��A��~�Em������YV����~�&J�`�$���lb��D-u+G�k�>�&(1���uJ��,���|�UV~1�)�7�)�1��N.Kh�����+K6������/*w�1i��4�=��GS��j��Mq������{�n<�ݠp�I���a���q�p����,ߢ��U�zn�k�'X�P"��J��b2�b':�j���ʣj'�F�V�0�~�n��j�}�����*�b�Ԣ�JH��K����I��%5>�,����Fz�*��U��N��E�\�y'��Yg�R^����P��[<k%�e�J�W����}��	v��}m.l�y[��'?3W�ۺ������G�Îi�(��n��o.��{Jh�@Iќ.o���Rc�F��%`�S��G��!zb��/z}��3!N?:UQ5� ���\Ow��e	�C/̸QYsag�l]H�R��d�iVϓ����
�*Z;��W����>,
uޞsu-~`Ǿ�}JW��w�)mξXι�Lᯢ+��an�Z$k�^�5�YH/Q��y�m�����@����_�9��~R(v�
c�_Q��D_1k�CM�*PY��.`�P �����b��)_��UUg+���پ/��8)�k�9�
����n��M߬a�O��G�r�W�}b�l��n�Q�\��X�R�5.�M�B���������̈VV���*�Vj�љ�Lw����M����m��}vu�:���`!P�Ǚ��#j%z=����:W���ǨYuf	9;����FC�;��4$Eq�geI���(0?
� ��vyHz�h�˦`�h�E<�:�,$O��d,`�?D�NU{�v���;�Oa���_q����6;r��� ~�b����d��o�S��OG���m�c�Wrx�%�5��ʗ]	����N=��{fe-��w�t�g���؂E�d�a�\V�L�ԅ�Ve!���
�|�L��nU)�/�y�Zl�ʤ���8���x�2ß�|w�0�F�×��8��� }ܖ�M@�nVe�^=X ��R;��-���%96�:��"��=�ƍy���h_�
��/�b\:V�ǩ��Æ��XJN!U��Pw�!��-R�?��w��6��ʃ�=}-F��6�j�jg��4����_4��nhJ�?�K�ȴ�뾸����Cu;H��U�>a �ڇ�PeԵ
Qڬ�;Mb�Ƣ�ۘӬ�f�u��z�MrAbF�����e�|�$]�&�~�$h�+k{e�/IXP&�<���}��W�V�/KS�q�1�?�Z� )���q=Ǐ�����q�%���ޏ�����	����{+%3����#�0D'ؔ� �P,��:n�o�D2<��=Ia3���y�N���-8]����L����']�����wİ�A�=�j��1��!}.m�3���M���Xt�?���-�&\�_SH��ȱ:��|J��F�����,�p���e�N�<����������EvL;���Y-��o��E��Gp&v"8��)��w�)�k�X�Ú�|p@��o%����0�����d*��4l�Io�v��l���|_ݣ._����|r9��2�ً�R�dw��6�U�^���͔�@��?}�����.l��N�*GQ0{L��Ǩ�'�R|y��rM0^���;�	���_j<����&����L���� ;*E� G}�s*d� i^�l,BZ�Kd�.L� 4�SE�VѤ�䌝�E��/�QD�wd�`�(Qײ�I���~%dT�՝�A��4���Ф=�. >eCmR\���T������\cL�
/��IL�� C?�Ex��
0[�����A,q�O��
�e��,`\�"���Ć8:�O.����i�&���R��&�d
zp�i�M�����9��JGo�q;s���ҩ_�Ǜ�hه�v��ʯViA� -o���;A���A�fvMM�]10��~4#)��J�(I��J ��?E�od<�­D����+��Nn?��Nw-�A$�k�[A�CpV 3/����uI��[~��~����>�?+�/^�l=��щ}c��m�dg*����R�yr_���oPp��F��:w� �ܑG�,����S��ݑ���N�����=s���9+��{Zf֒��b���\����{��z�U\��P���//��f�����GM���_���כ��ښm��*���L�b�{VZ��\!�袻�23��m�'�2,rrОԭ�&x G�}|��6�� ����J/4���6`�1`Nέ���_0r��p@��c��hc$UɓA*�:_a�JF�b��m����B�{b=�&6���l� \ɠ�����s� ��8�!.4���o�op��癎�}���� ��ϱ�Ms�8ke9�:�N�}B�y�ea֫���+opbQe��Ύ@��\=}�L>[���9��T��H����%�*����I9�d����T������֗�M�\�MΏ�x3b'4�3��%�H7wYXxY��ck���,�"�wH�*h�<K���vJ>{n��7��Eq8���yg�W��jb"�4�^P�ni�Fn�j�?�´�+���K�[�� �, 0�V�z�/�(&�Џ� mG��u<*g���'��d��8D;d��Ƹ*Q�25<�=P[���F���U8��X@q���h|#��l�k3��:ɟC[�?��<k��r�b�u���FW�_��]��9������vOK��C�t��s�i�k�u��䶭QTP!���"��tD"b@@z	��CTz�F�J�Ԉ�҃t�#E��&��K@�k��>g���u}?�L�'	ɜO��c�wS}lY'��X<��G���a�mڎ.Nd���ϕ|mH�BC�����gb�6g�ӡy�M�i@i������\%�@�i��o�nk)�����z�v���|���QC�	��z�h�� �M4/Zw8Q<��ωEry^wj7�#�G��7g<�kgBW�|�rMė~Gܑ��O��;ώ��$��ڧ$����'Ԧ]��Ի3��v�_�B�|_.ofq�N����9]���}�'.�+i]��ލ$���e��(_C�� �{ F�\E��,��E��u��0�%�wEv>ZkY�̨�y�2� /z�	�Y�x}���(�T��;��mU)���RSQ�M��ė��`�S8�5����"����h��m9��AS�?���q��ե�e&$5py��o{؟V��;4*��{�gft�yQb�C�����]��
��·�����W,�wgҋcǽtHFa���<ڻD
�����<�1DS}&�Ftkќ]Ր�8�t��o�6��	�Ѯ����T�=p�1>�jn�ĳ3������׭��x1�$����d���7b�إ'�`vر��H��|;��A�!6D�?=DMSb��gBy�b2�Hsr#x*�	;b	��D���LJ$wt��* }qĒtP�rv������ Yͱ�N�Mռ���B��]K�f�\���o���~��b�����٢H�Ⲉ6�ee�9;�GR��̒��ׁ-ȏ�5+e1��m������.�Ex�;�M$<@g@�e{ 'x ��;�-f������:KƑ���#�w£��"㾖�it��t}֬Tɱ>}�����ڔ��"���~l���8$>Q�,��g�5��n\�֓Qtx/���ą�Jk�Q=?U�&�\ߌ�U/+{⍗Y�uy?>���vY5�fv�Q�uƕR�[��ɡ�@KjK|L��<�	���X�b�9���
2# D�X����Q-<���a�~����N�����9���=�h�os��$'n���39�IwZN�C�9E��=m�����4r�& �{�z�I�zߘ3�]}TI%?��~�
�ՒC��9�~];meҤ7=��0v�+�n�}R_�!.hgϚME�X9ѥ�=��qf��E�#:8��p��Mr��:pK�L}/��Fȑ�tj!�oʾ�����S�/�ëM��ɴ`J�g)ß����Y��u�b`5�KD_E4��L��N`%ӌ�1�;4<�Ϸ�NJ{@�Ռm�D<'£;��	�8���x��1,�ʃ'�m�bA�����Ȓ����it���N� dq~�f@�Lw��S��� M­��0dYH��1!�ѯ�KM�y�[�]Y�5�ϋ�"�Q�I2]#����|A�h�O��?�`��c��Nn����$���K}��Qg�+}��:��s��h8�bD�Q>[|�a��q��	���8f��`[���
���:T<��jĺw�Nj��W���~����*���B^$����_��h��˥V�����/���6I�����l�P�C���]J֪�r�U3�C���J��\4X$�I#e�!���LD�,h��3v*�g�����ºU��6���D��p�$-�+	(�үܒ��l�>��J�;���AX���O�f�	�2��.pL���.��f�F�<c?�*��瑴;`?[�0��l@�Ij�.3D�����*�bM����A��4���p��T��e^*����o��ԫV��.}]�QڷJ��(A���Fռ"��Ё�h�*3�$��|����G�.u,G��Mvᬿ�Vw�=��v�=@��Vx%�5Ne�0��p�2P�ƶ�g��;��)	�.�9�E��v�/gJ.��L�.���Ý���eM����5
��~�)���өoO����tK��mY
$�C�� �f#�l�}���`��M8`�g}��FC�1Z�<�d�P�m�i9n�ģ�!>N����z�y0�h⩶�D/���r1�۱���s]d|�@>�f:Y�bd<��t#������hit���mF�{�'GGw�Ш(m������ma���/�V��p���ˋ�;[��S���n�i��f���r�Ԏ�ſRn�%-�ѥ��-��¶�֪p��M�ɾ��I�3w�+�TH�~b-w�԰Z��X��i�%�W4������������u���ghE!}�]��UV��b�L$>�o��7�ii��6����y)�������Y#[,E����ws�5�+�v�냈D�1��,�)�v�BXN�CuuPH����a�C���h�� ʢ	��s�Yq+"��4M|8����Ҳ���`����L$qȋ♋��R����'�h��}A3>�&~i��y@{�1���Qς��Y��A����l��^<�+������4~��"]�
9����po}�b�k��w2����b��v,}���N~�+VG9�3{���s�l�Yܴ��Cd�;��U���Q���y�X�3E��✖È��1�L%�Ę&и�"�wy��)zZo��_���KV=f�Kߧ?�Bv�9N\���1�
LW�%�	ۚ�~��1{T�A���Rw'5p��:yՋ�M;n|�y�]S7nv���"X�m��;��BN:��d�����};�"�Ҧ��29e&'�jJ�3�S�t��-�d�d#tp
��'\�
R��zl4,_yT�O�0�,�������9�$��X5bE��i/��̓�$Z�T��Q���u��>�"ש�wሓ������?m�J� }�����d|�ï�<S2��</�'�7�}r�:�gr�z>�$0��O93���N(q@�"��Y�<-���z2��F�RT��Vk�:���8�wX�K�	�@��7sT\��GFϝ�'7i.8i���De7�nt�ĉ�������\�'A�$��Lܰ��?�q�og,@��u0����:y�Re@-v��WeD�<�	Fr+�J�Lic��(����C��qJX\�ic��w���z��}(�C'�ܚ�Q�9ܖ�cn���X�dͻT��=��X9�&�[�]T%���fM���vt��ժ��k�Q����V�9��C��wnM`�0��^0ؕ�)����r |��*A�|��LVPU�\[�*�ى^2yH���I�&�(���a�*6�6	ֲi��i]�e�{���]q�do�R����|��
пt���P���Bݮ։��䝽+�跨��ӭ>(�%\ע��_jO}��)��7����������'�=>"N�7��>��K���RA�KqV �7Ȼ�@��e%�9��@ۼS��,$7g�-(�_{��H�a��p��b�ɋ�3�#FkZ�3
�UF�v�/� ��_�,Sj�9Ý��F#����3`^��T���/뫞�
;����k���h�}��0'��������������mk���	>�<"�N:�]�˒�.���%��G0b�~���;(�����>b/� ���Ř���%wg�P'��_��:Ǟ��%�J��%dڝ����/Fe�At:�|j���y�m�3F���"�g�~w*��/�%�bMw?[
�3]=�K���1JJ�LÜ�M��<t|��Ӌn��Z�]*�k� GZ���cX���Kq[�e�栄M��c[ĲZ�潬i�*�0g6.<B��#-��jWq_}"uMډ[Fn�Yct�{��q������1��ٽK�o2�k�nx�H��� ��� ,�Ǝ�Ⰳ�����!鿜.�d@b��� ��|�� ��Ƣ�b������Ǳ��t��*�[ͻ���vg�g�Hg�դ)"M�;�Q�����l�������[�'�	��Vdפ����^Su ��n�tD|��p'��5=���9ɵ*/Ú�Z�8a̰!���}��ѹ��|vl��-�N2��>��.�ǐ�w*���Z�}Iŵ��őS���0��/U�C������Y9�������۰�m��H-\%A���ȸ���p�Xaa�j\߃'��:��*�.u���p��I��J�W(�C=��+*F:	�@�/� ��+����7�3��������sp2 �  @B}������y\�>��QL�
�|�f�Iu�����o\[��{���dv7����>0�CPlu���J!3j��x�I����,��������:�>U��}��%ـdJ0���y�T�-ڏ�k��/�e�"�=�5�X�S�$>�ڹ ;D9��sv�t'��E�6���HZ6Z�.�zq�5U��x7�-���&������"�_o�����rv�T��@�Q�u�}�CR��$A;Ӑkc[���G>�U�<�syrѲ_R-�}���h����o"��_D`2OFNF0�KKTJ������ݨ.����� 5�d��v��S������0a֎��M;x��ܸ��	RT��c��2��H%�	BŚ}���mj�� O�x@x���qW{K7��`�2������a�,��d7��GN���n�c�nsa��Ǥ�wK����E�_�6t5c&�S]b�\���2�<o���ki`w"�B�tl�8KS����Xc-\�2b˳��j�m��":�ICZ���a#�q��-��%�D�P9��D�[O^-W�zt׎rg�_�������mb�D r�B1��K7y�:=�iH�Sѡ�&��Z�`&���`~�Is�ix�4<����xoi�Eio/�~��䄳�ƹ����[Ć�v��7J����������JT~�86*�s�J�b�$�)C�@j3��I����l���0��Ȕ~0E�u������>��.���Z�Ƽ�ߠ
�I��*Au�A�Jk1��۱o���l�(r�N��O��d� 0c�[�/�6n�:e���ay޸ ���z�ǥ%�0�>���E�?�K[��0��];�e��-u�R�К�CAug�,�}n��NF��ֲ�Ň����+޺ �0�����'b�o�Э4x-|wB�R�:��o�vY习���QB����ݥ� �_���XT$�Jwn�X�z
4W��������ƣ�/��-�?.�5�e��BsG��JXW5�u�U?�_�DNo'����N����>�$4_hΎ�H����<���?	�s"�����	��9H� ��uk�o�V8o�Pnj��ژkTVGq��������S�G���V��eOG�=D.���`+ ��B�7�ңy���vio�������!X�V�
�SOB�/F 6�`�ޗ}
o����p���q�7����$l�[��w��v�C�����mܱ�da��+���=T|sf���_���S��x��H�%$t6�;eꖓLZtz���Kg�&�M&����~�h�2Gy�MwQ�
���E�2�{t�)�52p��	�u�����=3�e���`�Zy
ԋ�,�\�\ڥ_�#�zy��b�W�@[�����\���o=n��5�mK��"�纼$i��'��H�RM�����#~N܁4W���y��=�8h'��vq�w�T��_&��+��}_��rYK;��y������sF���^@�lHGZ���4�	�z�;ë6i[ٔ�\���RM�|/t��f�S�a�[ox��h����(i��	v�Gn�$�ɩy�>sqc�R�]J���.�W�7�np�{��W�Le�`��}�>���)zȂ ��f�N2��g�4�" ���zV���&�W�3I�o�oړ����dub�?
�ꯀi7�Ky��>
ݙ�_�}���?r=�d��ä?
Yp�}"~� ���4��^[�,�8�a���D}�z�b8�i�}2��<E��:���`�5���Ł�­��:u-!4,[W�H$��k�߯X�#+"�%"�AK&�&��۫x�6v�p:�x����K�R#^�w#������pc;]�; E��bBK����%b��*f2�x,h���/�E��ڲ,�&����E轰L���n�M����.*��������n����p��/,�*�������\�o]:Eͨ��A�;Y�Մ��g��z�:����h��]�ڔ����Xh)]�Cq�O�9L��n��n|H�j7�Fؚ��um�n�� DOr��äT���/aI�m~ea�@;�f��0�p�F�dPAY{��oy�Fl A��A0�E�j�ǰ[x��E�
�g;��?�� [����lo�d])D�������a�X��mgfw<B���ʛY�s/!+���J08�`���4�1L,Y��<|���Rn9�Q�c�>�=dC������~��iA�V�����]I�Y���`���E�/��:��v�����X�'���u��R�󳱱g��&�8�g;n��h�խ��AV�R/�8.����7�aA��7�$�?�ó�"��`�e��4]O�?(7���z�/�&r!��:?�]uh��zH�WH����t##�WD��S�[� �VxM��8Q�>���-��h�����|���D�C8�{/��Ů��Z�<���f-��ʻ7��X�4�"�鯅���<-O+��^|�o��K8�0Ŵ}�pj	9	��~5ˌX]Z��z?�����B��W�q�g$��Vk�9|*gwۘ�z��ka#_j��{ ��U��5z�_\<�}�+@��צ����r�
��%9�f<�*Yz�Ғ�P*s\M�4x���p��.	=�q�����Rp�cf=g�H�]�c�(�����.�7��ڀ���L�N>ඓ\���L���f&y�r"�̨��V.�s���_<vH���G�%cD�%�\k&Ek�8�<�F�7\	8qI@Ɍ��+�wb���@�f�1�z��^N����Ia�:p2c��r��񅛱��!�[���г���#��w�	_?[��[iU畟�a��9p�o;�U6���v�%�fWm��d!v$+����&qxLK1n�f� ��a���x*(7�߮|m���[~KX��PR��|-К�X�x7�NLM��3������ݰ/�O��r%6��H�D-���y-%��Z!3�M?#a����<O���ڋ���+U�9F���V���i9�~����t�8<�����Gͮ�(���۟����ϵ���R�髬�[�q9��SIK�z^:	vg,��)���j�_c�x�B�#r�\7�Ma$Җ;���G_@�`m�wo.��ht��K�'d��� ��s5��f�N�á7Y�e���_�9�4�%t��B�[7�tw�m�83��	��9z1߲�4�ˤP��;��K��DzQ#��rE��vY紐��~��������>���9̍�m����?)���u�J���V�ٹG��o��ʩCm�h��uZ��5N@�ў��"'r"�	����~��q�u׊[��%��,hcsܓ���۩)�;q�%�;g{h����d��}�Աrj�;<��;rgH�`���-��)]=:��$7G���V�2v��y�̭l�=��߀4z�8�ɨ���V>�>��j��������	�5�5� 9����C�H�h�o��13;pi����X�"���Z�*�ٻY��c�E��޶��,��}��a�A9�V�AF�Y�1�)P`V�KM��9WI���Ⱦ!�gԹ��'����'�g��@��d@^E��#����ŭ��Wk�b
� '$�h�H��]�^�d���md-'�`��EM�~�`FR����17���v���Я}�vd��9Gz��� ���Ks����s��+6�
�,P�+YR=r���nKŎ���x���ի
�T��_+v{�FFB��pI�E햓juG�)|���� 
�N;!z0���a6�q��\��"���2���0��C�_�%y9_���]gۀ+�t8=��e��w�F7R�*TK3F�� #.�6 sFP'`F�����]{S��{�߬�ӔKF���㩄��:���U��3#���R�n���\:W��z�o.�U�J�[߽�Gqҕ���G�-.�r4�Ug��T�*�V�m�"���-��: d�-9=>7���{�~�հ�h2�f�<#S2�j����i�,� ��t�{ Ӿw�?�e�~f����wPn$���*�L�g!�<��tGYC�%["$lP+\{�G��kHX]fڍ2�nuy���A����k�m��n�tjB<N[�[Y[�$�3:,�w���L����W�5zF�§hsu���կ��wMq9�O�/u�z��N�_D4�H�!��9@�,r�g{ vVĮ��Y ���1�e�~�g�9��R� ��5�݈�8z����p��<iy��/���ߦ"p�챿l�1�BWߣ�݃����ǎ"^�V`��=�ם'E���o�3g5|l]��G�*J��,�q���A�z٘h[���˸�
���<�n�ȶ�gz4�u���}uU��~��m��� �|:���;�Hs�|�*�!��FL��Ig���<�_E�ִh��,|J��f�����]W�?a��?0� � M�v��:�We<��9>��/U�����}t�����|?5��ӻq�#��1P�B����W�����az����Á�=��``��_��چ�O��Xڽm9��=Z&=Ǡ|�)�CqųZn���K~G��A&�����Vf|�i3o9ߐB�>�440�4�eg�O�F���U��=q�ā�(
�7Dm�a�����c�?Ho�s�C�}�Ɲ��%♂	�P�=Ԓ���p�v-g$]Д���L���N��V���;�W���a�k�CVz�Z��`�3(�;�w���^�`��~j's�Mu����?�����d%,�R\{��x�K�F�6> ^G����qw��Ґ�i�L���6�h��q��{0R?vk�XZ�@C��H���h���@p��� �����o�53�b��%1����D�A���-�|T;���7�.�\fn��dm1x{��g:��|���}�h)�f��������f�V������0) K�sQ�����.w130z7�G���ժ ���Y��|v�Ҭ|j�D�:�<.EhH���ĊI��E��s�a*��5�5����1sY�9<�_+�2�Y<o�i՜�p1�@B�>b�29�ol�b�������jHw�!�;L�A�����s�$�%�Y���������ښ�?�.S����������M�xy��fE:�j}nw�&Ɖ����C�w��%�҉I�>>S~|E�,���mH��dv�P2���L�;$`kʼ՗���8A�#�{LL��QpH}@[������{P@w��������X���k3��]:?�Nj�N������=�
�`Y���KU\D�b��خ��|j�+d��@f'����/�>?�U ~!�R�f���c��D/"5iO/z1�<��7��"TF�n�yOM��5��!��,��?*lchnR�Fq�*Y���[�a�J��E�7��V�'�����P����� 6<<�r�� �8��w_а�c_�a����D"l�0?��s����%}�ܚ�$���rY��4	/ܱP���ǌ���H��;��Fۙ���.Ҁ�.�s]=�(5���G�]�M���<%i�rH��������u+�!�RN&��m���{����7q�)�\�6�Y�e�!�h�&];$x�&��H�YN�Cae�;Y�6�E�3'�wض	�9j�s�U6�7-�
Ӄ��Qv!Uy)l�R��"�G3�'�IƸ1$��҂��/��2ƺ{���y0�������������r��^�Q˻�}�� 6��xo�lu'���sg5��"D4���]m�c�6Y^�ц�ȏ?���oM��ז�4�&��:A���) =P	��GO=K�=�s�!�j�5ZYM ��寛�=�dJ.WE�\">,���Xh��!��"�6׻��F�SW�yK�`��e
�o���d+��=��^��o&��7�
�27��/N�i��d7:>�|��������� jLS�*��\?�]�@.~�c����	Y��UkL�22���/�ܾ��{�4�);E��a��m���ɥ72#��϶�zǍ���YWh)Px����z�BP_��I�RT��R:	H=IJ�O?Ƚ�j���"~������S���*�����NQ�з�ʻ*�)֐�9�����
/W�J}]f(��[�ǯ���Tl���g��m�X5��i�p��dY�6�|S��H<{E��S�B�������9��Fg�@Ksx��+���j�k����;���^E̍<}J��>eb=s$���S��z^��\��V���Y��D�����,Pu�7K��q+n���&\�=�r�i��m���Q"�:�{R��W���V���N�����)�I�:T~����D;+4]����l�Wʿ�"A�lv��z�����hDRu��/=�ʜ�nx�Ք��	'�����|)q�z9?�ğ���X���ӵ8z?��k8�x�����N
88��J[y;,�kw�׉I�/m��^��9�PȂ&.2��1|*�윕aZ�����E�\G�_�cZB�� �i�f�m4"_o+��g���9i��b�� �Z�7�BX�L+}�wo5��va$h��Yy����V��jZ��3/��ݡx��3l9|���?���$��K���gL�7�+ 4�}�ǳq��/�U6a�:o���8��?D�:.L �*�M����A�8l)�K1Y���¹�K���ѩ���O�ON�3��b�F^?il��4fm�n��#:]!�н���������/-��Y��K��z+ڀQ���Fh��j2-7�U��.�5`�|�|b�.kTn� �:�A�d�U�ya��b��e�t�/�H��V��;R�pa���
X��3�d�X�5��E���Y?�y�V:�K�s�x�w���݉*�DO��^���*�T�}�m�� 5�������S=�D��t�~6>�}N#�P��	�h-/�A���ޠ�Y)�ۙRR�\��!\�ӭ��N��v�H�҇��ؔ�۟�HK���-#�&ʽs��i�f�
ex���_3��UX	K�Hhc���Q�[H�I��`�Y:�-`�;��~�lc|��/ 4b9ZmW�Xّ�i���n�T�,�4�H#;G��\�F,����^E�鍢�HS���{d"$2�����{�{ R���#���BL*�"�c*��(DM3�$Dw�&_*ё���5�:"v)�� ՝���l��<�W���є���L�jT�5�� �#�=�w[���"��7�jV#�F��/D�"�#�<D���B:�=@�*�Jg��|b����.�A.�)'��qk����ZHH���!%`����k>����JF��h}>wk,lB�g����e}Q�ʯ�������M^f���DtK�r;E~ߙ5�O�:+�-ߪ��K|>��twty�L�O��j�ä���h*�erz^����|鈊e4Oݹͱ�e���n�������;�j� ט�pZ �W�2��Ҙ��_���8NeT�а�9vEM���q�����7:���
�����S8_�z���r�ɰ\�u��*ɨ���T��ҩ�Ů�s�	}�鿸;�;2<T��-�,k�a~����*�ߕEe"� �}<w�TΗ��EN~[60�<�q���ʳJ� ���5��-�T�������QNk�+���0�a��8�:�腙P�{*
a�2��Wa(r1t��8޳"r���#��|��G=Yo���?��`�-�3ݘ�CSנ��[�4&��U�-E�m������T�a�9�唘�Y�V�O��EE�·U���P���/R�ܪgc��͢Q�6o� �ݠ��D�>n/k�g"0za���O���s�u`r������Պ��E�'����O!W��|�+nGb�^��6-P�$R�6�ڗF�ZvNwT>8η������/|���%�@��pj:��.�y��NL�/=?򻡸�Z�g�x�Q�n7ͷ�����#��	�"�D*���py���d�r�>��O�=Cj,��7�{˽sF�mc�L�ZZλk<xY�v���i8s�<EU����/U��n��wL��c)`�<ޝ�O��(w���J�ur�����)�Q�l?�ڊ�����pp�6� �>�<��HL7��pZDF8�ogk�ڻ�H��P����o!z.��9�i��H��^N큼&�i#��ަ,��2Tt�<_��,1+���s�����JT��v��� ����2D�":t�Sk�z?�p����׀��$�TI��Yr�
i��ֳ�wm�@Ss���Hf�	^K�k|��<7�l�~p�U೫�~���h��n9]���R�1dF72�Ur��ыa};��{�`�6����Mj�P�v��P�'��~�3�ϙv '�#?�4�7��@�.a+�ϸb��u�������*?_�;��E���8��0�w�bhխuh#��h�Uf�X3)�Xj�[rA�P���s�������|S
W)�����=��[gs8oF��=������n9l�]��������j�s��z�l�k/�Je��5>^��w�]3⮎y�YP|�3�*��%���P1EYb:�;�V����r��"�%{��/��"�A��vZR ��	ZP�b�[���2�WD����7���ۛG,9V{p:*��y�Q�����Ɨ��\-x�Cu�'�����C~!�9i��V5��k�|��X
$�Wu����+4#"�k&a��_F�Ehk�,�GuT��sf)�������7��j2[�����'�v���
��n���u&߄��s�����o�k�#�����%�eL$d��1��<-�ߍ���U���q��= ����CF�3���$/#duy�/�����t���������`�oʟ�D�����*��{�/���k�{��G�-�=�,lkz8QYEQe�
L~��m,�[jJ�K�����M�jVV�K���ЎN}~���?LVs��`:^�'��r:�g�o��gJ�v'?�!�ȯP�@�	v���v�a�w#!j�L�<S�oA��I9�������I��7c�N��Q[�*Lq}̒L���r��Ox�O�?"9�D�c[\�BQ�+�:by�s6��_R;��*��wU��������G*`�6��t{Q���c
�Q�o�)�|�d��'�����Tf��-*����ܙ�<� ����*�'1[�;���X�«O��ܱ�Y���Ix�Kd����
z=�'�H��6V�9��6�ߥ=�2�o;�5�嚯S��&ҧةE����d��@������cz}\�%{ Ȱ���ؠ�/�O�Z�z����"4�Y=u�^�;#`����*F���)o�kF���������ǒ�N	qd��?G|����LN��ᣡ]	���z� ]�s��$-}a#l��E3h\��}���aoF
[Q�����t��#�$�V����,��LMm��{V+R�*ԕ@����|����8P�����d�Єz}����W���W�gW�����E�y������`�x��V���S�=��:)ʉ_5��������O�y �%��Sܡ:�[�"�ԅy��>��g팂ۗ)� Ϯ���@����:P��r���9��C�z�?$����Q���}Kr�䗵�S]^ �F����yH?������o�*�tG�U�-�m<�L��¹����/WX�=8g���[m.�A�'�H�:`ΟZ��=!?�|���k�]̒��\�r��~���,z��L�q�@���iF����$�pa)�1��G?t���Az|v��m�X/S�ŗqy>uJ%ғ��gF/it8[	�;����\[98,�ټ"&��woe��Ȁ�����zoh�yk7[R�_D�e���w�a�iD=S����_*���(�O~����S~��Sf$��HWD��qR|,U��s�Nv!��(Z�gF'����Uwc?��5ŗ���+
�(�����eWW���d���5,�vχF�h.u���LQ<�x�6�ؑ<p�+��퉮�e���Z�q�k�媺��R����Tdw��[�g���x��A�����fD�_�_���S�h�����	7��AԆJ=�k����+A�9�\&�8�-2Xu.RF�5�z'Ń�b#ǆ1�+>w�	!>a����5(��a��q��.3�q��N���}����ܽ�{����z,��Z�@k��/�S����o^�R���˿#]2�?��
�s�YD<�a�h��CY:�+-h�Ԉ&�JW�)�����7�
ݸBw���z}�7-1N�:�;�_����(�<��a���¯�JO�}JOFȏ��xq_�h/m�]�p��7��)s9����t<o^��S~!���5I����pr�i[�ë�l����hk�6�����[�����Ո��{����$;ͻ�. ss��Su���c��9=y����7�[��	N��i�.ү�~��8�p@���6?�a��I�5���\`���-ʢ7����<��\���(s,X,�O�4�����J#���P���Ǡr�Y���c��������ތ:�_&�L�EH��7�~�J�K6(4��&΀t-��ti}u���:-���pT���V���1���8�r��.~P�uK>�}��B���5R�p�=� �&N�`'Z��A�I=߽��kb�o+8B껞z�@U��
h��ݼ)�O���$E!jԳ�s���y��bUy�>��<A�d���a9�)��ij�J�e8O�/����8�L���t������J��7J���'�'�	���$RF�ͲL�Á1ǟ%}�6����`�I�'���d�t_h�@��h�-z��<FLEԗS�<��S�H�Z���R_�0�pb��0e�\/��8zƼ� R��a�{��W	�y����^�''��4�!�Ğ��k�T3��Ŋ3Q�+o�O�x��8h0�Y[��h��|�=�m�s{��=�)�=�ջ�-�����y����nة�	t��6��#�'��&�" ����,��߽��Ԛ�g�tw7����N��A�wBƼ�a����/t�Sh�&ԓ���mn�c�� oLj�|�g�tNT�U��ƲoHdi<{6�og�
���]6�mR��<@����}/ aļ	���Chb�s��r��$��
u'~-�\9-j��iu�t��Y2�păT���JO��Ǉ�!����<�f��;�a@���G���pJ��(g9i����y�[\��9�xU��(	7� a'@D,'�&)� �A�}�t�'3�3��RsA��g�}>CCxn�x�~M3����J_���la+t�E'l�F��q{���= ����sX����|W����(�?��aY]�֒Q�'�{��CC����>O��T�#�QQ�"��Ug�����޴����[��{7B{G�=7O+��u2�.׾��S�(�p�O�H�ό���sv׉�Rh��G'M���d��ҝ����Rn�eu~�Bjqe�'t��]��*~�+�Y=f��d_-����A_�/̧�P�.���O�o���J�0C��J�����Qw=�ws=�WM�}t>�W����m�H~��!�'Tv��-�C�����X�m��h��ZimB�[��5H>>���~�����Z�2��JXi��.�h�Z���r�/��"o}�:��x��������+����:O�Hm9Ū|ğ7���8'�|��艖�%R-12ml@7��_m2W�e?�+�U�v�Ҭ�-�ɪ�s�=ӐW���8�$i�ޯ�BB���KzI�q"B/ޖ�W:Ǹw�\:�e��O�+�̡���֯D��N_��0m>��ڍHI���T��a7=a
�>b#�<�9xDV8��Ҥ�/h���W�q�vRj���:����~6�);x�*��n׽��li���e�y!y�%N;G}P,:#��<�Q:Z|�)�r� O��9�kX�o�U���N�֩`۔5��:M����,4&l]!!*)+�kp؂��F|#zfN("K��̅����USQ?��%�1Oԟ�X��i���3G�!^X��<:�]m#Ek�CG)�98p���ZP�{�-sT����|i��lti�a�I,���.��fU��ߗQ�>�:2Ki���(M�/S�i�������X��UK�0��M���F�%+��*�TK�U27ls'�(���(y�����"��<���{._Z�����s�Ö^�у/�lq�R�ׅ���tW0�N�5wgFVr8wЍ/�|�y��|r���cj[��h�����pl��#�s���"F���j��1����f�k��6��
\����������>�2$��)��r��tEo�̊���Z��rl��%�,��/|���k�5Hތ��5�e*��%1��7n��*rC�v�x�v�O�dz,w-�ЩA^�i�Q�c4��,�]Jʱ:�0�}�(*�eB�)D�og�^��gD�}|O<��8��n΂=��r[;H�_�/^8pӣ�^+�j-��m�0f>,wf�\�UY�������X�]��r�21�\ ,��J�1�����9�D�)��g�P�7�S!�^yJ�81�2��u�)4�w/�TB�'���?q��T�k_�)�kȯ��W�7Cyz�[�tW|�/��\B@O�2@��Y"��� Qy�ۃ�)T}WkU��B�R�^��^���`�#�Y���i^r+�ћ�G���
�d�Z5�kF�L� K�2�$�<Q����҄n}�JVg>Ӎ��4T�)32��/]0���BY5^oH	q���%��A�Ò�|eDB|�'�<����wM_�)�('�1����-+W�}(Ƞw2$����řP������$���U�O���f��7�=�8�Q��g}p?��l�=#{Ϡ��2�׺:@�/&(a�[Tȍ�$��N;@�T�e)�XGn$@������]��Ҡgf��',�����S+B���?��@����▄�j�e���CҞ�`қ��]�{�,`$����E|�ǎ[Ló𱤉�@-�n:�`o7�L�_V�7�"���K�{�_��ӿyϟ��>�Îg!�*u&��{ .�2z6�~��������~�/喝]����,^����N��!To��P��sAz�kχ-1b�ͳ���;�$rG�;ysk�®���t��@F�\#d��,驰@+<(�u����y\��uW�[{��y��l�g�c������0HI�����^�)�L4sV�	R`z)�}�Jc�;���x�ÆӚ�����m���9Մ�i� ��9*��7���d���/h,Ӵ����XJ��MA�hU^��ml����K�*B1���;w5��\.)��x�yƭ���I(��f?>;�Ni����<�qr`�
�|㽦��b��)v���>���Z2���FÎ��'���b�� ٮW�;��.��l��6���9XÉ��K���OP�9��GT�V+��6��qŎ��Hɘ��G��/�S_x�U��\����\��� 4tP
�n�.D���řh׳��[V�ش)��3�S���{i[Ϟ�!�@����;I��\odu���Z�&�_b�5s�W�+�� �Y8�rcҰ���w�(�٣��E�T��,r� �����ؤ����{�5��k��� ���R"M@�X   -H��H�H�N$�(R�K�H��ޥz�HoI�� ��v��9����y��t�9��+���7)�YS�X�@��7p����a�����5񕬾���4W���?�d�:P�����y����?(n��%w�u�(�R��
w�dk/��[�<l�� ��,��F|�Mh�ҳ�V�K�����J��_X��l����5��^�]bf�+�#r��c���t-�8�;�s^�ɳ�28M��Nm��:��2?�.�1���'��_��֫<��'������_tSd��ۈ�Ӌ~<u�q�.�/�W:'C�/���4쵰Vq"�7=�������[l냛�pHj0��]��5���}_���,�~4X��(�=Tָ�#[ZO	`'�\��y��]���.��!}�%��I���"����A�T�|0L�D�C���>	n	��b�yP��Yy�^'7j3��;F(i%���(��=g7���O���O,��S<i8c����d�y��5�@{�s*�7h/b|��]�\N�$7�^:��"�6��m�{40�-��I�a��Ė�0D��	ȑ{&��Q&��N��lS���F1�ˬ�<�}AO%CE�1��?����KM�x�?[wag?��y���7�e����R�#Y��@�/ڷ+š�+űy��,�铴�#�J���I�ӊ?��������c2T�^z��7����J�z ��^O"��8�o���W7ٔ2x���^G�]��с�5�����7��M�PS��6h��τ��B�n�	I1�1��^�^��۠�*�߾�k_��qY������ �D��*���'�¯�lN ]�+��df�"�������L%�[ZaV�.p';&N�Qtqc�6.1ߏr^ �a'7�L�0Zҟ><}���(J��["Z+v��1�9���G��@]>W��*���{�?� �T$5bSX{�P9ඥn��q�%�f��@Ӑ��Gv�����{�|\���8�d�A����8���;d�������Y���M�j#����ɱ�LR�l�r�x�� �ju�/��3��ba�Z��P�-'�ٲ]�������A	��o�<�鼶A��g:��xQZPKT��fi'����0��iE���ԩﱞ�H�u3/7g��w6�l<��;�%Ꟶ�ͧ�}TQ�m�q��:/�C7
[=���������r�����S��"��������-74EQ6�6g��{�)���h�9���x˞7$^,
.~�u�ҳ��c��V�bP��zo� �vQ(��Ҽʫ�z����3�����j)/�R6�%��x�_,u���������l�W�%|en}�a�{�Q��>� B�&���(�:y��Ҽ����m��qf��'%[��h��(0�t��ٜb�p�0Z3��y�Yo�5wJS�&��8xo�k��������,�_�)�\8b/�����MA���xU]"{�a[�`~~��'k��{�ek�/ԣ��n�أ�}�p����*7�@$l���mVNd�[���G�	<[}��m��A��'N&zr�]��^�N!S���u�J��6������|g]���(�6�U�L\U�V͢h�c�|��a������k�br�qͣ�� ������r����s�6��B��˗q��
�3X�N��<�l�kݱ=E�cxّN��Wm=�!!�V�����S@�����:�A��E�SY��aåP�ϖ4����w>�����>�T�f�VaNJQ7hx�K�޸[��ӧ˔X� ��ϰ3�;�߆����mPa;����k�{�i�sj�<��Z5���%�T�K� Axch�;�X�@���,��<�"V�;�[���a�$1Q9�85�B£י�0�"��Esj�ݕ��p���9aK:�݂�\�"�5 �ؐx:�щN�/�y�F�m�aE�m4I��պ4�[�=����}��"�G�"#U�x9a8p*���S���l;����|O袁�倃��m���
����1�[���ބg,v�机�Xt.���{?��q�e%�ߐ���%�q`���.����J�W��U������%���-�.6A��e����|L����E�S<�,8t�oM�O��@ZK�8���1�6t$�<Q�~�1z�xT?K:LSK�Ƞ}5u9y��u˟��ZW���ͫ���i��Zׂ�<�&��~���T�J�IG�H��|`O��T�����,���`Y��U.��4G]��V�ޢ����e5Q�L!�A��f�������t0��c4��XyD��in�JkM'V��T�����U5��nR�>
i:�ɯe_8�q5!(�K6����a���t��ٳ)�Vb���6�#�%����͘�����:�wG�:P������ZMv�Ɵހ�tz�fXM��#�b��8�u٬�Z�������.�-���8T���m�dwbG|�JZK�Yu�#��7�?e�� �'L@�.���v$2�%�}�
Wp�}z�k�f�L�+A2H�����w"�MdI��&�&�4�I���#Se)F�ɴ��u�+��|�c��������*��"�אG�m�l���N�<V�tADx�'���.�e����̒4��ˎ�j�V���1W[KXg9�sOZ�ӎ"[3I�F!�G�-�~�������J�:2O|3?K(�~��]�F/�:��x���� o-3�TH��t�-H���{<�B=�ŷ��ӏ��ѳ�+�:l`ڵw}�Aa�e�f��|f}����Nx�)H`zf1O"��eZ��`�ß�!�h����T�~��h���i�}��ve`��֗b�&F}��Kv�W1��L�Z,���S�������׶A��0���^]�+�9z]�:�;��.�����[i����龑�p�X�D^Y�a��N���s�z,g{��*b^�j �77).&�g�XUztƄ+�n��@���"����iR!� ���҈��kq1(�鵿/��q0(ߠ�	@q������rl�RU���s1u�=/�)�W�P�w����	j`�|+��.$��?�]VQ�J�K��E����?���6��;��Y�8�+��m� D���TZ���M� f+2ӱ��<�!Ӭ��fO#�i��g�Ѭ�:�� ���'4h9�.[��$r%d_U^,��%3>��Z���XNƎ��Ⱥ�7�b�Tfw��cߖ�l�6(
�@g�VM��ν���M��u��f�y���,��(���5o�����X�����6�@$/�~�8�HW�Q,�I�B4'cp��5�m�k�,�(V�����f�������t�|�U���zF����m��j��e�����{p����/�nܻL�<��Wobǰ��S@L�H�w}��ݿe��Ԗ�����]�����x̑�J~��G�4 ��?�����MՖ��r�Uߔ�TJ�a�w�-L'BN���٨�U?(�N�eZ�b0�ʻt�7;�q�ek�����h��h��ݢ^��ΧQ�K�il�1���7}]r�I��y��{Y����u�+�� v�7�q���+u�bn�#w�����Ax����}���n!����O���"�!u�Q��&߄��GC��b��~�ub�>v���]ٷA�f
��6�5�;��p[d%���F�pku)����k����l��꭯�r,)'wHҘ���N�_i��*c-�@5�O�[eG� y�26�΅6��Ca���o�7 �?�7��x����j���eÕf�/t�c�A<>��u�_���m�HV@�5�04[*u��58�(�!9͠���!��������b����BA;.a�.�K��ܛ�����+���ׄ�����{�=^�q3��A����*?�8i��~���W���叺ش3�n����˲���"��,�eڗ�f|3���L��hFN~-�B�d �(��Y_�w���^(i�,���L�]��������\r��&��2$>k`/�Ѡ���ѩ��5�w�mAx� ���I<��ni�kJ�@��ۀ	+�#�fE��ڽڂvC?�/�'f�p�
��f��aq���?�9؁�#;�Ao���`���x]*��l5�:��ަ�o��:��Uh�a?�˿&���&&}m�w��li�E��W{��X\=�Ȫ��&��3O��q��,���Ll�hq�#��!g�(p�Z�C�A�:8:l�^;�<���~w&��7D�F�:�`�����}���������@����U͍j�.=�C)/'�y�WV��w�ʝ�a|��x螝�Ɖ%#�Tv�Sz���)[���纰Wn����+?^�/�e��l	�l������aˢ�?� ��X����@�o��%��L��_U�LC�*S�Ʈ�'�����vt��cÊd�A��m�^,�f�I�����a �0�ݷ?&u����:��ہp���ī鿣�$���ȐHhV�bOJk+l2��A���[�!/f�!W��
�Ve�������?�x�;�ԁK�Rw(�}_�>4K��&"����9P���)��Aq}�����wv6&�!P�A���̭����8=ʭ��x��Ê���$��4�}��� ͜t��YM�m�a
���>���"0_��z8x8zUcv�]��.Y2*�'w	8%����9�;{w� �K�����$�=�����6s7�4�4l|2��uj�ˏ�2��e�|�+��#$���#Jܪ��{U��RCI\�R��?(Lod⭅�ʧ��{_S�}�+��:��5���D��J��1ӓ�]=�ļ*{Qo[M[?y�S<��b��~��1��M�>���lbfj��B�� ���mE����'�¼K���������$���@�g��H�(�c��3&��|�TCK	�dތ��"���'u��4'��ݭ�3O�#�^CGg��6S#���yԫ�������u�Y�%NK\ke�Um�_�a��8Ǹ���6��iu�"���L�*I)c��Էd�mЗ1'ꨕ%2U8`h�0�
�v�xGN�ޛ�č�˱�J���2Ď dsڽK�ы����o�-���Y*���wpT���xt�w��ר>Q���!,��q����^���(�1N�i!-�<�ۼ����R��zN3���S�K����	��"��FZ�嘳A��Ҟc�*���g��^�V��H���ǟZfNኌT����2�Ã�=@8�;@VC��) �z�^�X���@GjH�����I1O�\~��j'��q09�UH&����WLh�+���f�ik���!N*��h�8�(�5+*p0<�Qaպ)�\Y΄��ퟎ#��YjG不��p�Uqr���Tn�=̐nG�O�2rz�A�P�K��of�a��������F��uS 7*h#3v&%3��������I7�gא��u��n#RZĵrb�쳐���c>���a�wQ�od�[p�3�ثC�N��b��-aP�\��|�L.#P�\�X��@��,<\S��Q��.� ��FĒp'���	,p~�B�,��HL���mv��ۉ���4�[��U�(��(W�F�EbɉK�����tH�\��_hǇ���(n+�ܛ��J�LU[<�3lS�z�I~Zp��H���kI���y�eÎ=��ӌ�@�����1<�#�����q߯��?B���9 �`�ud��y�P\ږ~jü�1F�����c7�7t\����$b꜉�t� ��-�C�t� �f����������3��T� 8*���
"x�[{ܐ%j���U��/C`�>]�-?X�h/�od�)\P\5U6u�M���WF����t�{5��--��
��N��7@�����`�sdڴ[%8���xE�M?@2��^[����R�-ѓ�(�I�3�p�å��<�A?DX��� ���Ԟ�y�v��>;�|��ߪ2�!G�~��9ܤ"�����o�0p�x�H��5�t	�s~�6yc�~�i=R�7p�&�z���Z�*��þC_�ޥ[.̑Y�UL��%jν�ԳO��͛�,�kX}q<�kQ/Ż��;F~h�׵�몔�˖��B��tgq����yIȜ�c��;�w���*6��h{ۤI�L8�^�gXe��o����EU.�u�x���ʦKU�u��ُ�\_ŗ��Y�v��z6����b$�j�.�	X�5�'���Y�1�^�+���aw��c��bҲ��,\�f�\��F�a�~=D�&��z�*�*���b�s607<?��ϥ�+2ދm��=�CA���>�4����j7���O��	��$D��,�,v�HƩ��i���ݬ:�~jT�|�)=�V^��3V�;*!���!� /�������/k3�a��#l�Ӻ�͝�g��Z�FҎ�P��j��y�Z�vT���4kP����E>z�p�׏髇Fa1Y9�'R��j��^�k�j�탗��!:�W���2�z�\A��%�B���#qr��X�`��+�+�V]�\Y�+s��x�X���g���:�t�:��t�{�"!{�8!� q�(�_~U�S��rHk\fS�`h7>�����.<��&�U)f>A��)G�b�Hۍ�ݔ�L��[���e%�1cP�s:ړ��%�v]Є�����5��Xr_0��9�q��L������K*F�1*N�!�4���S��3(�j���<�y���1�h0�veNG�J��E��֬_�`�G/�3�
S?��T�jѬx�x9Lۂ��	!�?EvIA��:c�K������_%���Pi���>"o	f��3Ɲ���{V�	�z>h2HM���r���7��٩ΓV�|�͂�V>&#�����+�'~�B���N�m�b�]��D��e,��u�詈�O"��1V�r�2R��EO ���H�DP"�� ga�������u3�wQ��;[5s��p���H�o���O]���>$�Qg��ֽz�@��z6�|p������W����p��·}���E^�s���� �6�UѭO�c������ƺq��;����G��v��-�뢕ߛ�Vm
�@�Jz�^��o��޵��_5�>���c��Jf#z�1�_�����E�q�9_kn�}��Ծ�U�\x"V$EFP� jc��_���=����#�ȅi0�;r̤:[�czH�� �/�����e��R�P�n���e͝��\�&K��@a��#@(�:�+������a� �W�s����gJ�l\�;��a�+��R&~˷�|ޣ���E�§��(�K���T�LŅ��rP��Z����6""m6��Ik��_~�m�F��Jm_PdE&���X����J����9g�Q�D��XlOY^�͘�bSf�{�Kǀ�M{>-��@�_C��B����t�!�5:�Wَ[%w��	�j����\���⏐U���̟���(�9�f5���27�ܤ�7����]�%�]Y`�M� ��]�;:�oҘ��Z=u蛟�tA%�UH�MA���U��Se�]8?i���a�s9o��ajr��OO��ax�K�wѪKU~L��[l�_��$����N��G�f*� 5IF�h�����1�����uf}��4]���tѕQ�33J���KG3$���؝<\C4b��Vgk����-���=I���o��S������N������dX��8]L�nխl�P����z,?�8�5Z�����WK��)`�y���f�⫦4���⸙�D�f�5�'YBz�3���"�3S�"��U3�@�ܸ/����>w
;��Ā?��{x�F�[��%S3���5��y�zFą�8�#�4��OW��@<�I�4p�&�k��S|_=	hs��fN�Ĕ��A��-+�gk��(��<�VWTW�βz���3Xa�e�tLůg>�R���̿b�ڪ�0�+��%�mU�f�S������
z�:�qZoA����z	:�T�*1¹�ƿHN�}�g��2 ���F��⁸��ր;g��^�4�A}�Ӛ�|}t�J��\�I��i=m"P�~�����b�\����_�,�Z��B
eFg6~�AmM-�����n�3b|˛��VW��ސ�4|�����7�����fG�����!�tj>d�UQJ��k#;��s%��ő���<"�|�D�����D~l���I�1���i
E�$���eY���E9�Ӹ'V��f�TjMzG�"u_?M��9Ih&`q��6q½�*|��� Q^>�5�h�3�J��L���g�5e�axh��Y�W�������V�X�G-ok�1z�B	'��rZQX�R��_I�%"W�w5Ց��(��W{���;�z��^�`�vT��}�p!������+"݅8؋vy	������~�zο��3��=��p1@���0P�_C0D�ಠ�X����;�?�ı��ۡ�!eԍ=C.�>�U�"���@�=�ar]�u�¢�ǦE��_�Ū� �e���z��=d�>w�W�� c��T��j�n��c;'�o�!�:yO�X���D6b���������J�]%�۬Oґd���}Pй�Of(�v�#t�)�����I�j���;gT�Ν��re���ѡo�~�'���n��v� �Y�e�Z�Q�@�"B J�$ғQ���-ƾ⯳ճ��*������b�4"M�A��G�bP�{K��������x�=��݁6��j�~N�Q��"�u�G������I�̷���^1�-��R�o��)	9�@KF��o�<�"��}Ͼ���k~ϛ�Ɋ�fv&���c�����t�̀uL�Z�(u�>'�mP�����N��fE'Zg�ӷU�/fuZ�Yj��w����� ;�5�71z�?=ϵUsm���Q=Tgy/Bz6�}��h��t�� �zEn�����������'�3�4���o-�3��W��_�M�)���(�3?n�;�@c.�m���b�����N���D$�mq��ȧ��bʱ��v���RN�`�f	2�f�''��[�ε&�G�n!���O+>��7�ƔFJ��T����0�
��X^D����ɓq��#'�*����O��Ҷ��p���\����dⁿ�i[L��Ӷ�Ò�(Dd��$�y,餫q����Z��#DO+4�|�s�o"C�^�b�DC����H3t6U�e�{�,���4���������S�|���O�����6Cv�Y(�>XDt�9����H�����m譃E��
�`��׎ ���Ym�S� Ȩ���x��h3�J�"�#�_�)�X�{���o� 1��~3�:����K�$��z�U
pGl��F\H9�[�����1�y��tHô�8���览����tnn��\''�7���H�]F>�m_���87����
2mu���UE[�����a����ځԨs\]���CF�ߘ��E%��](�x4���!�n�\YW��;Q��j��l�h�A���}�y��N�K��<��a&�'�c.�$A[��)��CLN~�b�f�*<�ڍ��m�$s?qh���1	$`;���ڔ�Z�B׍/	!ʠ˧} [%�h$] ��ĳ�<�sC`�\����-��
�K^7vX>�;��dX�^��U�M�f�zn�o�F(LYx2����f1KkY�F��W�����.�A�[2r�n�����\�8+?g�6�H[�RCRgh�u��{(�bg�`KE��������gRǫ���Gp�(���zyHz���V���M56��zu2OٽNqT/b�z5����a��8�>���^?K���ŵ�ϯ+3IH��Oy��]!�A��lB3e�h_�(� ��-�|�����Z�(�d���9����1�&ɏ�>w{���{I6K�Z	��+�f����sp߭8�	c����@`V+:FK�&C�mͬ�+k���.`be|���4-`V�@�ɬCd�XՕ8J�E�>�I~�<�F�3`���nR R��լ0��f��v�x�:Ѧ;�V甧+�'}'���U� /���8l��g��%�ٙ�~<_�+љ;i�Y�,�8u��/P���j��߲�e~Z:�X�^ ���ƪ���z��C��5�W� Y-r��w���%��:����ŧE����B�kP����O�����x�g7�2�
}vj��-=j�b
�w�{��J��,���
�VT_��GP�n6�l�R2�gi�L)~�r�!�Nx��B�v�S��b��H���"�gd��̋�"NYށ�pX^4�жo&��R�Gz��L���3��;V$%��֪�)y�������O���KK���I�ǅQ��z��q���1�8���4.�Z=dM�=i��N5 �?�&{�� Oʴ�N���6���x���7�tQ�0��9i`�C�H�km�ʮ���e�\��_��r���?�H���bt��J���7J��q��gC��x��}���S`F�m6���[���E�dix�:6>�6�ǻ�% �k3�iˑ�rC�<g��ӊ��yǨ�9;��"H\�V���y����;��dg�ٗtC���x}r/(D�Sh�����S�G�%<�nR�_F4��Ԙ�L��_���͟�$ �۪��r��ų����D�Zv"X�'.z����}���uz�J�_�~a\��0���z{����V��,=+�Ħ6�q/d�d?lm���x�NA��\��[��~
�T	E�(��\�Q�s��!'����RL��m�)yg�K�����,O�O�3Pr9��ߓ�AY􇔤f~5c�p32�ų���8��C�e�y�ޫ�#)3蕜��˂�r�p��t��?���"��|h��|�!�Ev�PrYCL���������q��7�p~b����	v�w
!�de��0_ì	�9��gL��bo�-Weƭ��
EN4�y�����W�de�-?Z�g�3�2T��j�����iS9�����x�h�=��_���n=t��e��=��AVM�e�ަ�����J5�p����L������͝�C�N�1<��th�2���g"w諯��"���f\��N.����Bыޘ<Ε��~5m|4�ù��u��t͈vډ5�x�fB1>bKө׫٘X�|6ו�?�\lV~�v��`�����{3����H1������_{ǃ�m���sj%[a��p
�e���n�W�36
<ֿs�Sx��Z;{�#�1��^���#��Pf �6s��u�;��i�lZ���o��{�j��~����,"�=���f�f��鳏��Ma�/����e��ƅ��o���P���V�f�ı�π�4[��D۔q�-xf^c$��6��M��l��FMV�Ը�|kF`��=��z+��C�k�KVN8�Y��)����A�zA(�9��Ox��|�5��L;U��`�5���o�E^�©+�=4g�NWLU�tW��K��/ݵ�32*���-y�9� �C�� ����tUU�6�riEh��R������x�8u���;r\1��~��x�W��t�_e��cFJ�y+
�	�)��4I�#f�9�������?0�����X&XRf�_;�W��T޸m��
rmb�CcE������wJ�������q	_��������[�~����$U�� �-j���*C����s�5�#>��UԸ베��q���S���{���^�h��nm�� �㰌~ҽHn���Xn���-Ӭ�z���,%	��\�h�y~�Eb'�'�-��F���d6r�f5��ż&���DV��Y�Vf_9ۃ��QZ�`GRo�������:I�����Q��WI�>)�O��i���+;i�;������M�G$��A�NR1�>��5�+? <q���@��w�a{����kj�_ۧon��&��Z� W|=����<�2�b�%g����b�K�b��ϗ��n-[o�A�L��/��5���t����^�B���;{u|��"�/�]��^<ߔ�5�;����ZS�[�����J��f�?��Da��"�隍XXULp50[���]��{��y�n�^���\�t�|�5����(P��ft�I�.t��p����	;��ujP=Ë1���$���Z{,�C����b=>���f��QYA:<����G�;�'�1q�����D�M��ך,7L�8��y��?j���$�!��T����BW�n۠���	C�N{}��𝭟�uQ�n&�J�ipF|wu�N��}<��fC��; Fs�=ʤI?����u-����>Lnk��>��~������Q���+Ӱ�wlA+x�Ў������3T�Z}�r�Y��Y�0��&�rS%�.�Y2��x5��G~ekOr��������j�xe�< *�O���rW�rЎ���;��D���V��V���6誓J�d`��$#�x5�g�XM�l��ٓ���n0�d.�S����V��/�.}Ÿ׊>Ύ�z�_~���O�����C�ֵXV���x[V��))oc`�%a^A�w3`�O��+X&��}+�x��Zzt6E��fT@I)���7�O&U"��j�[�lr:]�X����zm{�&���t�Q�l/����<�N��y��ͯl_yf;e=1���$�,�3��ü�ݿ�FD�
��a��Y5�����d�ǡ@�����us������i�ʙ�2dYCt�e�Ͽuno�n��KS!��)�5ÌH����h^!���%������^��$��>�c���E�[1�P�~��]�w<rx守i�	W��������\��.����y*r�mĳ�HQ�')|o0���m���$�Mʰ߃ܲ�D� �k�:Q4c�^�c�'=(���R\q1C*K7c�8�FP|{��L��~�=�b�t����,�o���c�k�\�YO���8�:/�_�R��P8uj3��~�F�z���Ǳ�]��� ΫGa��+Qn�7a����2��*.���~���7������l<��^��PͲ��'��O����t'�{��3H�ZA�a#����ih�L:Ej�q��fF��x��-n���>����Hr�1��6��u��t�PJgM�R+��l�bK�J\�Jf���1�o��rtT$8-\��=�����6��d���/\�%�+TH����r�yIUT2������p~|gqך3KW�@���i��?�8���Т��/��'������7(��t����+�6{r_>/���W}�h;�/����U,Qܘ�k7�����2&�F���	��#��3)s��qh��6���e:���t��0�w�Y�t��ڀ��Gm�K۠��ɭr��t��Ȇ�����
���J\������S���ߍT�n���,�:Z�\�x�d�UQ�M�d<R�e��0���i�8_	7���#�_�gl���vL�e��;p=I8����A:B�Dųf]�|&jD`z]��H�0-��OJ�0��~�!T�z+.=��y奉Z��g������>Xk�M
7I3��ICX�ZNWF����!��_��ت����� Y���2J7�eˀ45@N�n���2��>4[�B��O���i��پJ�b�2��M]1�t���6l,����-҇��s�Rd�h'�k'���Z;�$�ȏ�����걍���+������/����_8�{�\�D���s�t,uU�=��x	��*��Y��3v׬/���5�������W6���<�[,?i6�9�k?�?���V.#����؆��0��K�[�:�QP�=��ƞ�tO�RSy�ӄ`b�J��L���tn�K�noN�B2�Wr�Y���	6*J�ם�p��-�o�����m'�h-�{��Y7��9b$���#��|i.|}3�u~�!Y=>�W���|��6-$�ޖU	���.+Ÿ{q@������QԵ"���,,��ũ�aNwW��EX�!1��P$4z�#�7!�b�`��@��KWHۥ�`~���?yD ѕ�A/m��寙A���]�O��	��^�v��F�Ya�x����u8a$�1j��\�l�v�6�ΰ
b,�4ˊ�0�
70�5{��s���َ4~2��6�^��z$�`��%�ۀ����	��ݙmr����,�Q�j�Z��K;˗0y�0�4�:���u���@>�l��.�P�O��/��p[��/�:��'�0pO�j����B[9Ƿ�G*�5g���i\i4d��Dl` M�}кd(=�c�9`,[#K��U� }p!j�nu���׽���~��sk�0�����(�~R] -�)���@�[=�o�J�_Q��L1�-cf�B�8MhY�7'�GE8�D��V�-�@�H�WDF�A�Sb �)BkPμ�����l�!�։(D0�ђ�"��حh��oV������K�Q�Jc��p_� ֢	a�����ojV�q^Qeu�<u�"�~&0�g�-R��27�w��0)��#�k��M���濾JK�ҟ��e3'I�V��T��n1���2�yO~��W����C��ݸ!��f��$l7;��6�Lڣ{q/u��^?�� l-��T��i�r���k)SM%A�-�y	ct���M,�����J8)8�����[���vZ����j�!5�x���-���M���v��thCR�b�\�p!���4�z2)[�{�N��j�)O������z\��5��6���H��̎���H��֥Dߓ�jZ���H}�:��W����sk�.e�d�\�~����g�xi��/�Ľ���.�����1��*��(�XAE��tZ�i����)Y�v�6���wm�hFRǈ��q�U&���,� B�H���b������y�q�<\Y����a��YjGL�D�� 7��N�*$�����;�����bUs����V�A��;l����r�@��쳔�S�G܏+5�V�NZ�Oj��QpL�rP	��*5�~��Hx���v������;��z�����Y����KMX��Rub�.)����q�ty�$��e�'�Ç[
�|,��'/1�;3�Ι�^￥�cV�!yQ7=|���NH������yq��E*s�#ɇ���ۼ)��Mǯs���雑���/���>l�g�J�ե+7g�:q�:��)m���f�0n�'|zb���O����Jq�ʺ_��>��b*KX���>d�Z3j� 2
���
�s&n|�	��z����r��=���+TD��y�\������z�����:C������ª@jfFft�N'����;��xg8�Ҫi�;[3���LI�¯�Yi��؃tY�D�&.���\]��si[���\��Ii��<�XJ.�r6�i�Ο<�fU�S�F|�{U�ÿ�]�blĵ����s�j�!f������d�.:��mVo>{X����;�dW!�Č2���Ro��xM�ا{U.-�l�Y�AnV���+�f /玽��lÎ���PiӰ,,~�5�Պ�%� ���+�s�������]sK��W�WH��W�^D�I1h,��S���qAc��P�i�o��g����� ��̗�n��ʩ̷�qM�vl�ʜ����������X���|`�]�ZP��pg��=Z��=�$(>��l�7���Q��>��m�*Ġ�d5Y�/���?�b��\�����-z���YW��O9F��4Pj��1IҾF�2)�W�����)t�k�yaamR�|�
�(�G�m��I�7R�ٯI��3-���2�AA)�V�Vn�Gw��8]r�_�R�h�fkUK�x��Uutji�+�Ĺ��Mlv/n��|'�4>�2k���}V&&j��%s�u՝���،4��>�uzXKF${��]~`��@�4MJ��@�����Qt�oro��9��r��C����$��^H,�i.���>o�
3�T�	}DZQ�n^#N.C.ݔ�$�*Q��Kb���	h!䟚�O����'.�bN#7���#��eG�)
�g��V��tD+*���?��������O��x\��M���~\p`p˥�0� ]�:��'��J������t����e��ݯVK�"�	�^u�j���>o�`�镯!~#��ȳ9�"Of���ڟ�E��˖�1��B��4�҄9�`=7�U��.�R��v�s�f&a��z>0��-U�z0�2u�n)W�*M6ȕJ��Le7�5�����{>w�S�@�'/lƸ��c�	J�7·�v�?�U{����٫t���x��Az��2jS��ff��|�E��L3�c�d�=n�ы��
�z&e
������ɫ�6��.���c��W�A� ����
tF<(�jy�
BN�ϐ�4����OY ��I���N|e���F��H
?ޔi}j&����F�bM�����F��bΛ��d�>����b�k����eڴқ�>L-�nUg0��������[�2�T���t�>����+#��>�W�i�� vq
 ��Y�Y����<���倄bӲ�.�����궊��~_~�������6���2�������i�XK�[7�-�/_n��o {c��h����
��p:Y'0d!?��ǉ�^�jG���/i���ɑ�R"�K�1��~��*�_|��w�OjQa�P���fO�Iϙ��:c�5p��/⾽yq?L.?y:WL�%��V��Ì�(U�;I���" ��|�/���E
	k�Bt!����G��Pfs���"]��?�ٛK���eh���t�@��^͟hM3�Z�Qm�%�ӄ�P j��e�\%�v��у�0҃��^��)[�\D�0���H�WsO�(O�9���o(8*8侄�]��L(��=��#qD�`f�5�w
��(���!�g�o�I��	���'C�n��as���ҳL�g�%�p�A��-���:�D��V��:p=n�/���\WH���ڥ.6-nA~k~���K��~���PJ��)J�=j���O��Z�:�٠5�}��t�����~�(��KXcUplWQ�Z���?꓀��՚ܑ��� ] V�����|L��J~I�ѥ袤�^�E�
��Q/�����W���>�>W�~պ�ŬE��c2W��?�œ����vԻx���*����yZ+��z>��t����4~�o�X-h����7b�����^�VՒȝ:P���C��0w�sp�Q��]����G�*���p�ӏA���CU��E��S,l��%cuG�T��=|��u���5�4���g��'s�[��=W'�E�4f�'���7l���8�W��_3�,�Q1��6hϫ�d��&�� fҷQts���H���'����)8���7q��Z:51��^iN�_��4n��A!鴒}��6c��ll�S�����i\�'�/��DJ��P����F��o�ZM�µ+�9ga���T�f�Ş.Z�%��-F�T,��������F2��q��!x�[��-�$��湤���5�w���61�se�D<^r�߰<��B��u5��}��	KC�N�$2�<^�F��X�=�dbBE���^^�:`5Q�W:��C�������<��> ��;�>^�H�}Z�!��r�-^<=��剈+a+�o�'��Q(�V��������=3�+�ëi���;FHO)<c
.a�0�o�@�I|9�%�Z:g��x�笂f��.��ʝE}���&�ԃl�%m��a<�q��Q�ai%�#��i�C{��u"�u峿�R�R�����aMl[�Q��X! 5�HQ����JB��RUD:����D��J�I'�t�(U�.A)RE�$!��P�s�i��w�w���?�	ɞ={���[����kϭ��馤�m�pHh�K�`VC��yz�|�(D�c�@.�[N%�0g"������q*-`؜�$ot'2�_IҺ���;�gM�沁�Xuel���o^�ۜ`u�@��jUưS�k��A�����G%O_�FR����iߜa��g��a2�U�CDL5��n��l��u^���gĊ�E P`%�YSRwbٺ[�@Y<*���/x���ʧ��=����S6k�=>�y�cR�?�O�a#��vP5!������+�-�����0�����ϟq�R%&ꂜ�A�w�(W����Dת����*Pݻb��N��S�'�l֪�>-*���o=H�8��Ɔ�S\.J�U_�w�n�����b�\]5ˇ���N�M[��.�e�L�-n
YҮ�w���ic�z�:���^���s�>L�1��q���R��;��]y{_��U�g,v������OV�^��E���2�˶�
)8�'	I0���5�L���"g������6��4����(�!�!R�<ف8�	-Rh�_�YC�D�	��~�_q匢˞$K���H�S_?U&�N3�wW��_:xe�uzA��>}O����I���|��؏Ͽ���{:��$ibqi��؟�--�GF���&�9�0u��r�1���d?'V���?�.�)w�>�-O<�H�n�t'�|�����_>�y�r�ِ��1u���� º�<�Nrb��B����W���IG)I�t���/�Ą��z��ten��˱�1�+^�p������Ѣ[(_y�����).��O����k���I;=L�l^l/h0�D���BZ�x��[�d�lQ/�Zq�k[���������Ď�U�6	�=��m]=o��jI���~������S�~R�z�x�'ћ�A-I@���u�T_kP=�W�~� s8m[[�A�q���R�5$��� ������v/q)��=|�=|��<�1��Z��C�>"�Ֆ՘bA�����N��A�z�C_�Dl�ǿ	f��=��f%����.��Q9�"�{��p7�_�)�?�����k%���&�3�0�΁|�=:�
�GM8��Z�h�Є�Oь'F�
�dn7��g9$�����t�#��G��g�ʿJŬ0�h'q��ɤ⎂l��!J��س)+�ō� ���s�N�Q�`6:�B���H �͖|�g7�� N�Y�@{�YQ��yVt>���<dQ�2����]�K��<�+I���{�{�8�6��y8�Y�ԝ�l�IU�}߷ͷF��dWw�c�59���<K��a\��H�[9�V�xr|Y�S���L3�JQ~��z�T���V�.�'06z�:0M�~�&L�p�)��(�����w�4u�&�~�ײ����P��;J�BǷ�H;�`L���>�� ��Vt�V��X�w������c6%ίC2"r�"h$p��ha�s��/�w6��Z�"�Rݶ���,T��aoq���iM�o��,�N&���="Q0w��p��$j��Ӱ����E�=�!�]��O����'�8�҅��?�O���F���"h>a�|�u$���XS��=��{������-jړ+;�
�����K���1ﻃ�H�� �7���;�4�y�c]�x޸�f ��/�a��Z���r�v��]��p��K�xJ����G �!m���Ц�c�HoR�#���Gە��Cwqxf,��0~�Ts�6eO�⾇῅��:���O��Ph��J_V�ϝ�ne<O����F�~m��f�؝�Fh�4�4��R.�TS
�3S�w�e����}l�*�5W�0�]M�X�,�%������P=��ĲnJuH#���),�G��/�@�E�|z��]|������� ���YƤ=�qy�����Q�A?��I�~���V�7n���D
5��j�5�	ͥ~ų~�� 6�N�rx���g� 9GC��L�3�ְ�Kme��k+/��&�0�Q=�� �C��y���ӻOe�f��j���ؚ��۬��C=���^ut)n���lHGc���ϝ� }Hk��oFZ:��L`쭁-	�? �����_iI�=~%ϛ�)A���;A����%��e.�;)���s+�[�8�;�,K8����F�U)V1K}� �U|�2% �+v��(ArUb&w~d�^�!��Q���8��Ŗ�J��0�拨.���z�e-
�IN 5u��]g�@��]Y=i#�|�����L�kE�5)[=�cL��ƺ}Z���l�����[ ��L��|�A,�o������"��w>��v�BJkg�	�j�T%~9)�R�$r��(���z˥Xʨ�m��͆�}�C#ǳ���)}V� �2J����wi"l�����À�u�AR�߇��/S�@�t8��m�Tj�j����Od%��
(��r�J���Ц�Of&�z�����@��V,�#�Ag�z����`�8��&�!,�*���E"�h�H�5���{~M��P�|9�R��6�:UL�-�ΞzD�i�j4a�:&�J��J�C��
�<��s���������%�H�3��ri�]���m����$�{DSFN��y�/�:j����{4�։�"YiC��k^��p�xU ���w����a��ǀ�G\6�1�̮6�fL���zZ���g\M�vM�o<6�(�`�b�<&x����0��y(�6�K��Y��l�JD���9R�-t�eˬ�ˌ:H�v�3���=�����ٶ:��u��i�on�u�i9ڗl�4�|Nzv�)T�q��Vz����*��`(�vϽw�𤿵,��0m$s)��i�:�E�
����E���]�}�k�����j��5~9g��န���g��h?}�=v+��e�˳�2E�f5���>����!o�d�z�E�e�Ǻ�a��Y��Ӝ���o�{A������zx ���(],���$�|LSŊ�X���-�Я�௾�ϧe,�>ǔv��%�sk�@�{{�g�W>E7�*��9�{�R*����g���えw;���^g��pѵ-ȷDj�e��YՔd��sr�����-r�[���������
��2὘HcYT}��{���dV�O��t�T�*�j;�{}!:�K���]�]�A��g����t�8���I�6��?K�CK�����P�a�����O~W�]s��O1�:gXL/��寈 Ɂ��Y����Qg1�"�U���t�Z6�kz�mba�o����,iv��ê�"V�Nrf'��� ��R8`g��n��i<_��5Q{�9��X���	b���m��� ̤�� �ւTA�mP�@�-��8�6OpM�0��7�]e�����ei���@���|Br���㱉��������2	\͑$<b�t'�I�n�H+Y�K܋jfGKn�k�w�#�?�~�IO��R|���,cK�ޙ�6��<�#�iP���(��+Ǟ@Y~a�xJbo���oh2P2�ެ����\��w�������[�>N�0�� �ŏ�\� ��b*��t����01Χ*��j���c�>��P��f] Փh1Z����<�׳x�շ����؞M%���\E�f��w�����}��@��%1�A�5Ӱ��k�7O��:a���gٝ�b؟ڎ?E$�J��$�f��J]�"P�� à3�L��N3�'2|f�m���J��Cp���	=��޹F�J8��VC;���r�e��Z�|�}E\.��F��B�g�+�T��A�W��ۜmDbl-$1�՚�:�&�)d�!%����&�,- �\�򩁟�,!��l1���&3�vC���( �1e@C���>��H����\<xv�ΣTG�dJ����I� =�L��V����n�@}~.~�'<�ޙ{=��Rg���&mgn�k������m�Woh�Qu��m��oN/�[�T����o�+pA�ߴ�8p=�S��i�4Tǵ��[�M����m����ₚ�zAO>�߷���?1W���4�5��M�ˁ�1*d��{ I�ǡ��D�vOJŲx>#A������M7�2WP\�Tw7�a�9.��h�*mPv�����Jw�D����㒏8�aN��:����IW�ʑ�>z-���E{�&�K������ק�8.�(�9%9wAiC���(+�j>1\�Љ�y8s5��6Əm@�_rKt��m����\ �����1�c�y}�j+	\h��0TI4i#(� ʍ��y���U�w��[�Y�H��7�:�څ�1�C��gy�<ևS��g�L�d<�3�;�-+�j��߷2�~�'m����{j�-T��N�eR��>�Z�}���D#�������Ы��5�P��f���,P�����9�W\ƆeNi�D�;ߤ�G��?���ܢ��p�?�;C��ע�L�PT�R��hu�l�c_g�sɡ#���<
�s/���1����𽑔,1��_˰}Ћ�� ��@}�6�V!�k�MY�Go#�f2��S��$<��������O�T�[�*\e4�l"}�'ǆ9g�|�'{����ky?����j�G�;xgL)xN�MU/�N�3�Au�N�ݭ<cj�zxl\.j��K�	�:����RF��j#�JZ��:�Ȃ������S�T�}m5��k���ax'�B?���#�^���N�2՟�	!�hEZ�K?��R����u��}u؝c�H���F��>m:��q#����=i�sa�žVyU4�9)c�w}:)�:���|сuc��u(.�E�� E�4>��-�i��&MƖse?c�)4v�A�}Æ}��J���Ѱ����F������jųj�C9o��!�WYN�J�G����Z<��e�ڃ��/�Z?+4��p�gi�h�^�Q�B_���^ms�����h�k�݃���հ A>E��ca�ʵ�6���\��ZZE?��E@�6���/�^�rE��y~��1	�ٺ}��6�����|c����Â���!';�Ύ*��?��bԪP�=��jL��Nf��N���	Y�����n��vһCr���mXy�D�6iK�ýW?�b\�/8��(�i� 4ۅs$G7U�ɚ"ǂπ������P	H@�|NHg�Ǯ`��~�fhk�u$fM�<mOyۈ)� �F]�C9����}X���D��wذ�ÁS��H���P�Yl������KC��f�B���0� g>��^&����]���t�,SZ\��B�4]	��'����>5#���Ĭ(�}E�T��a\z���,N<�H�9f�5^;�?�	NKCdQp0��<���6�.N�E�h@������?`�[�s�5�?��ȕ�~�若���fꐑ�����7g�iT���%�ŕ���I��IһzF]L��|�F�G�e�[	���6�SP��!�F�S�J*r���+I�oRJ�l�����r��6���h��ݽ5QA�~�Oٖ)�f]����8,��rbB�5^��{�{_f�j���tپ�����ˑ�
��l%���1�_��6^E�\�i<���D�n>����i��o���xHx�wFy�?��wb|�޷���(5"�I�n��_&���$\L�3h��
�ȉW~(~Ć�� C�Rφ5�?��k^|��+�6�t�*�4�Z�3>��Gݽ�!�ƺ���Pk���{�7ݚ �$�ii����A�;D�wr;����/䁯���'���%�i�AhN�?jL �ւ�W���\._�9�5�%j��d)�{Ѭ����$�1D*G�#��Ã��/\K���)�����KK� ��3�k\vB#�tL[�����|؞̎��{��[!J��[��K�����3��Z����/�����83�g�l�f^���f�
�ذuDqs��>ږ�=:4h_'��b���R��j(�D�KF0�8�@3��^�� �hl[��y��#��'`���ǣ��.'�lǆ�	����
{̃�aD��)��0KT�U��Ӻd�7�ڋ�ڋ�c+�^��GM�E�ŝ�l7��)lX�Z#�	�����dj�`RG��7)9esĽ����,��7|���iFA�̊���+�r���M���G�߀�;>�wg� �N�<�഻�����=�d���gb�M"a��.�P�;;�:_�P|�W���G��J58R��r��}��Zq��=�ip\�)߻�v��F��'s���"hv�e�(��!�I.�~m֮��fm*2j��q�ֵm���a=x�>��r��hj[�VoX��������^�Cw:�c�^U[�#�]���!�l({�Dm߷��>q��ϥ��B����!���BY�<+�a�ߣ��0����s>H�#~�2�[���d	�7�eӋ�m�S�<�|F
�C���q���_]�A\�ġ���p"�Sr3<t��:�'o%f�|���/� D=��X�N)�獏'�9'\c<���TkG	��󟐶}�����Mr��!��*�0R0��5�<��![���?�[�qP�ֳy͹ђ����z����.�Tf����6u�w1���h.�ܖ.�T�������t����k�ѷ��K���y��GstQ�~g���q�����[���v�k6�մ���B����+���O����-?��f��e2�j�!��3�-���%DtMbA�k\JC SnA��y�"eX���)8E� J{ٍK�
���Ro�7��H����������n�$�-~'�><9�^�_�[r[�k)�f;̔��&>86H�����+�/��K�����:z���5����k��q/����sowg��پ&���p��)e1�x�4ChH������]vB` k�=�l��v��ޚ������I�VB^���ϭ�Ѡ`�����i^� �1�̐.�ۂW�BohgO����0�Sz��K�ۅ[�I����q�U��oR��O��\�2�u���>���<t��/��a�������j�Xf���L�������AAc"�9^D�-�7�w�o�2�C�~��^jʗ��/��w+Cf[C	.�-������˔#m��5]
�k͞P��ʫfy�WR<�n`��R�%���1��|��_�^Y�L"3��b����,p$ �j@e��}�f?��|'f\�8����0��ʨ����D�W���9,\�h�E�iD���t��QXu��k#i/a����a8`%�t<{�_��I�v��;��O=�Z �N�-(�f=����ԥx���C���F��Q#�u�=��}?�aXG"�q��0�v�eH�y����<v��g�2\˶�
%s���r�8�Z��6�8̎��5�6��TQwh������b4�*��i7�l����o:�j͗lA=3=`��u}W��]�p)m�����i	���\g�i�Ú����Vս�syd�0%_~N�u���Vq:�s^Jב�-F�߷5����tP�v�@i|�J��AJk�����|�,��0fU���\������/l���E������V���.��dX��{d�mӄ_2a���v��Q��E^<oh:�hj8ܧ����!RM<�xw}|�E�▱��k�._��N$�2������_+�
��v���k���b-���e��\gB�v}�M��Z\P�ƶ,sI�G���H/�}N�l���^gS�ǹ�S���$ګ��+���=3G��??�����V�<uV��77slx����辠�f��܊�W��!���Ǟn�/	��������X�ȃ���WX�Ň ,��U,��E+F����	�͊�3��6��g�m�f���|�sx�o�s�7�L����y������}����#��̇~d�2�'r����P__<��)�:^}+���E%��0��\��"8�MǼBp�W��T=-]��K�f��7�Cp�Uᆁ����C��M�5(Ne�l�
�Ճ�Ğ6ć`���Ү�����|�s$�
�	[����"RG�3��ԓ}�h��="�KX ��'U9�B$@Ɇu�c׋�e�bH$��1�m?:���1���0�"�x��L7��߂��zfD��Y��`���Ө�=��;�꬞��2'�c�7��q)�e��f����uV�p�_T-�����Ə#1G�W���ao�2��pӓlX���S��ԫ
4}�	�w8V��$	[��;�8]�]o�v�#�f�Uv{����d�?Hڎ�,�����$f��y��J_��}5��G�O������x��짱޼�$�"�k+@ ��໹�\�Ϊ@��l�jP�\�/��u�L:P3n��H0�P}x��q��Ah5�C-���̚��u���Ӄ���:����q]��]w�9Y�G�Ê *���K���E���+o���a4��q�Û�����Z �)-���w"@�w�x;y��W�e�E9�"ir�/�ǃ�]�h?������b��Ҧf�
E,��ֱRJ����$��
�m=	�S�S�.,��ix�'�;Vg���T8o{R�<�$PI��\3蓔��oi�ua���_��ĝ}v���&S@T�m�H�UBK$��y8hyyA���m��"�ڥ�d�!e'Xri��+JLc��N��N?;�r�3�O�6�j�%��3T��j����}ņ��ʌF嫆��V��������Se�X������N��h�Z`�������#�~7���]X���`�M�d�h��r��a���-)@��?��c�+q�A��g�9]tej�g�>xhx��Ne*�!Kc�a�f�� � �ku�k7�n�M�G��i>B>�7N�1�� Arǌ,�q]Q�܉/EL��Oc�������Œ)Q�	�돡��W#��0���`$�t�C��?�O�J<<��������:���Ӂ�ڋ@ �l��4U7-t�ci�a���������&��͗���0�ډ��X�����+��j	
��Z祊B1���܍�$�Jt;��/lX�F����X��mU�U�ת�Ϛ;�#;.�P�(�}�T��!pt7X��^τ�I�F|�vέ\.Byq-�:
�'�lQ�Q�����@��b&1]@�Xi@�k�唲̀���.Rz�l�0��6?dn6��6%0"���[%z$Ur'��L��"��wXB:�6w�$;��� �d��{�"�S����/�.1WJ|�w|A��/,r������XON��X�ĸk�
>��f�]q�w�&Ϩ�7m�[��)  ��\�<�v�]
�b��jJ��4Mv��Fb	_��;�ҹ������|܏�W�u��4Y��6� R�tm��Jr,��5�
��l7@ڋ��%�11db�C�,-wr���px_��w�Y���/���/u�8p�a��{uh�,AY�#�O�����'�q�LT~֓�:�tv��c��ո%�E���ܶk���~ђ�ߛ�6�؂��\ƕ�V�T��A�������gR�Q�M���;��\�����ڇ r��H"�8m��N�Ȳ�bt��֒3jt�O����K�t4���C&��n-IB����3��:�ʰS�6,57�WA���ZB�`�pJ1�T���+"�"�5��J��Bl�AR:��2� ��ӣf��RepP:��f���?��a��S���_��Rb�/�}����;��螷
�	��'�����{��A���R�z����YG�'ξ�d*ϡ��c������^ိ4�x}v;��P�wH��}# �~�X_��ʱa�{Q�1F,.�\�vxy���yj/�b��1�ʆ)�яU��\�bhfx��-�D%���.���d��,�{ӑu�3 i�b�rJ=�W�c��-Mzn��s��'�>J��EL5�
�eFO$$�Oԟ�������Y��:��W�b6(�<�V!i��Lj�Yʸls)�Q�[#�^�؅��T6ΌH�$���!{�A��L�����o�4��ٿ��� ����w�3��oy����O���0)u��\�Q�БgSȘ��czomK�>P���)��ճ��g�����U�5o��m�A��[�:~?�B,����鱉f,Q؛���v���u^��.��d�P'��LS�ib�q{>�}zSsv���+�6�D�����"�u��|F��������@'�̻�B�Ѓg`�攴��tV�8g�� �&�kn��5a�c�`�fbX6i�T�Qғħ�7��_�&��{����
�#�����U��
�1��B$��1:�pR��	���Ǚ(�[��JG��i��%7���>q��A�c�04��3�a�!s�?�f-��,��$���C3t(*X��V2a�`�,���񍱞y��BM�|`�8vD�o�?N�o��b�@���[�tu��6��D�+�z�"�z����~+Lb��7/@L�� #��t��p�_���� ��װ��]��T"���㜟H�z�fo]��=3M �#X��IM�]j�.��q�@'\z&�T&i�Ϗ�a{�/��O�}���ˬs�G\����i��Fk�Sɛ�@ri)��[@�ڧ.�e�<\�#��Ge��5�#� p��7y+���H�7���p9Ne ��͍9��)�=��=��J�f�qsZ�׸�hP[p��/�Z���+桴�GW&��Ѕn���킾?����Y[�X�6"�6����65��� �(�ȯ�������!|�k�<tO�N���*��ʹ�Ѩ��<�Em�h/"P��mwfw�����'hq���+�u�A�'QB�*(n2��=���t�w�[zdb�L��ݗ����t�Wfy��6�P�<���1�9��_�_՟^==��=Q��T����s{6qӹ/QbC�X���T.�0�sFZ�mfȹ�_����8�o�wtӡ�v����{Z\	I���މ���0y�뮲��(���G�j���A���bQE�j
l6^���r.�%�Oֽ�qt�������0);;�l�!��X�����ͷ��PX�]
���"�����gP��şfUE��0�D�e�2~� �f����Ĺ��J6`��P�Q�<�q%{"�4�a%3�`�0l��W�������b�*R�6�� �ܥ�g�@����{�2��@h^�bk����9�laȲo�,{[h�g���;���́R}�!l l��/ac�IƝQM��	"+����\�|u��>+�68�+'kr
����8�_��2��U1��!�R}��䯙64t�,b�3��A��*Jc�92o�K�m��k׿0J]w~��bV��}@`����@9�&�˓��A�;��J{��͏Ė68�;^�?��l�	�jL��]T?TWt����4���Qர1�.�&���[�Y$�PTaN=���,KSD�U��T��LncB��T�'��1��0�uKK�M��&��ˉъ8�ㆣ���J4�7�82l[���A���<��3�����zh?���ސ����1Ȓ�m��!��Z�a� ��K{��f |���4�Q�OQDnG�g�D�B���)V�1�(%<��F�}#����������8�W��.j�5��8�g2�,�A�$~��I���C^�D�BG��݌[�FO�֜C�Q��-��&�3�����s��N�'w��h��)�o4R�[��_��^=�N%������?��b�w����yO�)��Glت	wz�rt��Jb�2���e����7l8��nL,v���)T1��Ӵ�x���sŽ���#G6�0�t��B&��ߚ�A}��9��|T[95�ݧ�sS������w���م�zl������E��)��O��U�]�B���r�SOCr�5��'�:b���Nm{&��Y�4����)!C�/�+�$�o�a�SB±a�fAA8�������V�
�5ԇ0���� x��ԍځԳ�WÃ��6K��<�g��w�ւ�*-�������4I��t���͸l/COib#����y����!���~k=kmH��F�~ω�c��I.-���Q��I2}:<w�
��z�dZFʗpܚd�?'v�1�렼��
[�"��f�O.2�*��8EB>��b��(̗$?K��w嶛ε�&F)\�'Ǎ.
�M�] �E6L�G���8�%����8>W6���ˆ��ˑF�g��1h��M:̓5�X3��f�����l~�	hf���k��,��%^G�G<����G"6���:ZR�뺵����6��(uOk�[5|�:ﶄ�B�i~6����>?�ž7�
@�c ��b 2��JD_�6KD��b���TO	��+<4& CS��_/-��>���!ؖIe�����b;��<�S��,�rC�������ߖ`���|U��'ݻ��Ĭi����|�@����Vf˰�5�J��;�~�5-�	��
U��܊�
#p�8LṒ[b��S+2������,G����f��|�43�.N��m�{1?�l�V>,�!k䪾�K;0w}��[l�_fEL��UK8�ʫ��~\u��x��؅w��ޤ�;&��6�Q���kD�Ol���4��Yڴ?��X���W�\��m`h������+$�k4e�άs)�~��p2|�%���w�~_^���~I��j�Q3����B�i���| e��ԏxnl��S[ݜt�O�Ӯ{"k�{r��}M�z�eGG��۟���P/.�s��P�(Ȝ��[���{�3q"+i��t�"��H#V-�k5��;K��Y�s��\��!H(T���
l�zN�i�S�$�|�"u�E�fVZ�A��~4��J�;r?�Df��r��\e��9��dbz��� lH�*�����`�����,��&I~���Υ�*[�����ް+��-{��w����G�#c#R�^�ċ}&�o"��'���H�Ӈ�g]�ˆu�zI\kbZ�a���ZM�'m��H�l"g]���ŨTA�������d7�������N�ǹ�\U���=e�үBrF��]J��M�K�Ⱦ,_w���g�
f+o9�X�8^yǛ���|/��!��m�A*��Fj�id"��=��T$�a��,��Vd��9��J��t⡀�h�֜�W���"�_�9�(O#	i�̘��Ĝ�֬��e�|����爋8���i�oyr����F�	���ؤV��w���w!��Q4�ٜ��X��,�����oc�����sڲ95�2��7�9����Q�5�f�>�^�0�怾������u�/4e�apV��-�K?�0-S�L� �Nv�ێE��}�����!n�Gغ��bF�.k����̶��ҍ�7� Ǟo�~ԟ�g�D�Es7o�ި/(IxwJ�HSD���hw��ұ�?�fS�HN�%�񽊸l�>���sX�;?�k�ZZF�e�JV�4�x��� �;�ְ�x�8�""����x�����"��s���׻X�i�&J�o'ua^̬�O�3$,���f ��C�4P� �W`��B��B��av�����Ec٣z��6L�PB�����m�a��7�ζK�uz��ܗ��<ˏf���)�H´g��Ð�ɸ�1A��D�˜�,<���Ko��~��^E!��*��hո�6��h9��h[C��b�P[eӫ����=V�0�xt�1p�gD�h)�>瑯��E��6����D�}bia�����D�w�y[�FX�e|óW��1|��>S�$���o��&���;�AZZGل�[K�J���S����tlH�%���_���<\	4�	���Z~�$|��Z
�kTUZx�.��Y��f�!�>'|P�&�������l�ޕax���2
����n�iS$N�fR`�4�/d�'7���Z��yB�qɢH�n���C��S)u',փԭz4tL��W�^�1�k���&e��O��v��ܽT;rJ��鐜��gK�&��D�DX�FtӶ�Pg���X���-���-�"s����BS[8��lg�v*����ď��`��p��������x9�N���nL��G��J ��&�E>�� � �5_��R�T�R^�'PO����Z�X�d�U���&�/���՞vcԕwˁ����g�޸w�4vCK�ڻoSuv��WM�_����Pg�s21��0W�'�����³���ذ��;�VxZx<�~F�g���&U�㧊ng�f�n4ɧ�����X�����F�HV�&9�d�E%L)lY���;��H�7���*`��}��UE��v$F�^�wm���s�MC3���C���ORٰs�����}�V�+��yi�q$Xu�Z�bu��Sn��ё+�s_O�+{ȣjr�k>s��5�IqX投����O%�m�0pv;{�N�}�<l)]�BDG�G�[��$�Ojf��6G~VA
��}��4�[�ȱ��5�T=R�[W�A|��n[S��=u��k�g�#h��S��/4?|e�G羐ZB#����.:!*1�X�.$4�A3r�V�if�H�?d��-��J�E�A���/�f���|��a%u����3�h����������������������V�c��&6,���z���;K���aE�#۷&�޷�aCbl]�_�.���Hm�$���ߕhΝk7��Q[h�ùR�KO%���!ɠ/��j���K��t��4M�B��+)������"fy�T��Vww��և�Q,�pz�Ӣs����y.7��Nr�Q�5�@� !�w݈R��@%�<�D��4!�VM��ʍ��uA�6F�J�I,z�YG����o�r?�p[�M��A��K�r�
�f��V�+Q�nΧ��<���D/l�m t[�HC@C�l�����R����/������'�O��B�؏�5/|��&\�G6���{�=����XH~��{e㙾��m�/4?x�fʴs�����{Cz��O����M=�v{F��ͥ��ǒG?��V���ݔ��88Y3B
�n�?PK   VH�X���P  `@     jsons/user_defined.json�[o۸ǿ��-�Tx���gw�m.H������FGre�AQ����vn�iKm���#?�4���ߐC�_���3?<.�z���>���|5����	N�̗i]u><�g��~v\e˼(g�(������>C��i�ҕŢ*�S_oF+K����`�s?�Ym)e��4 �G�p�$S	�a���视L��U�l�n�S�E��!^�+D�ֈ�8C�P��4C=�.���1����SuX�;2ˋ�"���/�by7�糩�|TNa�
�*�,��B�E���iY��Ф�$�ZT9؃n��y^��4�B��1�ψHJWߠF>����Z� Mm���r��?ï���$./"��.��4����__��곸>k����$������Ш������,*.�⸥8�����i�-��:��[j˨��j���*R��ߊ�xӶ���x�і�N��Q�8�-�rpz~u7Ǵ-����\��M4a�{��7F�O���M^e�@�+��&��u1i�+��bq�o�+���q�^ڤWv���x�M~e�x<��L�$Xv���x��M�eǘ<�OT�	�����9���%�cW�AmKh���Iw0�����q�Ķ�]�x�;�m�������_�Z���"�S�_��߭ӛ�����^�7y~2,��`��d�qֽ����d�I?�������f`�];���:Ymڵ��D�����������+U��W�|�,o2���E�6���YQ'�v�\��u3p�V��b��ޖ���Qy7{lQ�<_��<��ǲ�\�L���zbm��-�d��L�3�W0ÑC��N���SY�I�ħH+IQ`T1Ǳ�^lRpv����mJw��[:�I��u��Yw�W/���������}9��7�	��f�V�j�ASh�rJ�	�oR��dN�U�|7�|��-�M��0M�C�J�8�,���(3V.8�L����6�ލ���V���1�&Z�޼v꺖/�H�8I����/��׷e�w�2li����4�R�5� h�UcnF͍�.޶�,`�z��]����������1p��_��f��k�j-a؆���qI2R��ɄH��$����������������������������������������������������H-+[|�{a͈�2P���i�<R��L)��_��NX ��6�"�Dipy��Ti��i��$��ɿ	V�]��2�{S��'e�cliJ�O����������j�����R/�(��ܐRY�i�2D�`�
k�RL �Q�z�������SX��i�N�S��?�3����H	ɹ�� � h�!\�)V��`�+mR��Y�ʈ&ۜ���6^��aT'D*BFDKp~�W'bw`�:\�z.ojy�W�wq��k��#؍3�e��ٲ~�*�Ldptk��O�zp����e��m�Z;�
-i$�Y�L�%	�Y}d�j��:��h���N��:J`����9�Jp-�����G�=�(�\#g$�B�Ӈ㒻�hx&�Z୳�I4��;�/� ##HG��jv�A�����]������Q	匩=؁4�鷳ɛ�k3T�G���K��j��̎�?�3��h���fİ�aRr_7Β��Mƕ�(�0����tt~��6#����Û��IJ���Q�*n�	<��[����<0}��Yxku�<��䈃S"�E��<O�~�|N�ƈv���x�e0Gs��&�	%�)3����KgNkd+0�Y��=�HЌXEKX�?<����D�k�۰��#�����H�`������(>J��7nց�'m���[�9=h���r��A���l����MZk�A���׿PK
   VH�X`C���  D�                   cirkitFile.jsonPK
   |G�X�v��f �� /               images/153184b0-233d-45e0-a203-5756afb39f29.jpgPK
   �D�XYY5dl It /             O} images/1f408b97-f73f-448b-bb6a-3763ceb62f06.pngPK
   SH�Xo�>��q  �q  /              � images/2cd737db-51bc-41eb-8762-f3273c40eae5.pngPK
   SH�X����+  J  /             \ images/5644ca41-1cf6-484a-bb07-c2f9a6f5b19b.pngPK
   SH�X��p� �� /             �l images/7e81f6ad-0912-4ff6-bfc6-e58bb7840941.pngPK
   SH�XN�v4	� m� /             �1 images/91e5cd07-2a88-4b0d-9128-72e2f992e16c.pngPK
   SH�X?S��� 2� /             8�	 images/99226213-8268-43da-ade8-d9d07cfcec9f.pngPK
   SH�X$�8�l  �  /             � images/aa130aff-16e6-4627-9689-819d55b5861f.pngPK
   SH�X6e�b�  �  /             �� images/c0cd0a79-4e96-4647-8bb3-400a2b193618.pngPK
   SH�X~��a� ٮ /             �� images/dc707dc6-8489-41bb-a5bc-77a0670f90d6.pngPK
   �D�X�]B��  �  /             a� images/e79c4949-80e3-4485-be48-c961657b0025.pngPK
   |G�XEm��O �� /             f� images/f99a6fc2-4a50-4dfe-be0a-52d397e863dc.jpgPK
   VH�X���P  `@               � jsons/user_defined.jsonPK      �  O&   
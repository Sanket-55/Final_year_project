PK   �N�X�)��E  D    cirkitFile.json�]����W�/w�Z���o���@v����1`w�׺���Fc����~d��J�)��@���Y],�?�A�?N��_�V���}�����r����[���S2��͗����kw�v��c����q�j��n����-��v��������0��P�'F�RߒɋWc/C��%-*�B��*�Ru!dS5�W��M�L]3���5��)��#ф�%Q���-�ZhK�D�d�a%+�W$-�Ӥ�V��тZ�Ko�	m�T�j4�j�&�5Ka����pzL���Z5N	V��(�Jl����K�
y;��:Ž�p����.kcY���e!���-uSغ&΋�q�
-G�,p�˄���4�ܛ2(I��hSxI-���T�
#��Ԝ9�f�х�6Lͨ6[��Jiq�6D���⠹�Z�`U�41�j�X?pb��Qj�U-0UkD�%�#��9=R�h�`��H�S:	h�<~�P��"C�ko Ƒ�&*�L�T��9���j��5�dc��R�(=�,�j�����yʑ�c�<�H���W6ʹ`Ĳ����s]XFP
ͼ䴤e�{Y�)�T3*b�2b�.�lxU0iX!L^v�$�\;��M�� �$e��jN�TsJ)f�V��:_�����5̫0���6��T3�ͩq�$�Z@��50��������AX Qs�� �"D�)���5�\`�Qs�X������Ӷ=lbb'vzf�y��Kiq���	ߦ����S�&0ƃ�:5��v1��-��F���U��(`�#y�� Um���̍�b���+@�r�߀F-������Sh�"jN�/�Q��e1�,bP�i���A�
�jN[�������<�2��?�2&9��d f�0U��
pk��
�w侂O��0�j�Z#w�L�!^T�����Z&�4��$����P	���
��n�8�=��\�3Lad�K�Le�D�wd��.4��K�/և�N�t�EYd��#��ZYh&��n�7�"��u��lԵ�-KcplZ�*�k^bش𕍫f����8o0lZ [�42�6�I�#�.)Np<�4���sh�<*�e��y�0�y؈,���Vpf9G�򠘙�@�J�猣}���U7�y�L�D�<������ް0HB�Cpٍ�l����YhM���ͨFYt]�q.��h�B�Hl��f:�l
�X�Y��#M^f��.yq�|�y/�[<�]h��<v�9���44�a�.Z�Д\�e�E�B�t�Ah���RM��w�����
4�u~Շ���*�TS��֗h��,�R.g 4�t~��f�ί��L��5��9��B30�c3�lJ�12�"<�I�e�E�B�&��4r^7@s��74-q>h�0��@��@�1��q��/��f����Y.��?�KYX.�b�B�x.���s��/"�����Eg�b�p�yP�	�y�K�����/�`��4�i�< �yP��e��yP���A1˃b��,�Y�<(�yP��g2%��A1��bp����8��x.e��\.������T��\.N$p����b ��\\
�����ދ���\��rq&��x.g8���rq&��x.g8���ru��?��Eԁ�x.Q��\D8���rQ���\D/8���rq��x.� 8���r:>M���7��������&��󵿿�[��׷���j]����+��S�J�f�9q��$R5�r!S3n�N�f�����15cz[�j��uS3&K�l3Ћ�X'��1���64��I &�&!Q�xL՘��,	2`�E�5f'QZy�8�,Q5��D��0U'?"����W-�nj�\��9:@��a�똚1��z����15'���8��	�@4��	��s2j{�S�Z�K��+Q��0��7o��ڿ[�.�[�c�� ��s����Q =��<�C� ���9�c� H/�� ��,�@��gx�/ ҃�+"�#}V�g��`�j�X�:�Nv	���Y	����K����n�x+B~'�
��"`��� 7�`�ؘ�Y	�#4� ��� ����W<�}[<�}�^��Y�Og@cO�,ACx	Б��p��a�<��;�����=�k�?����{
z���.�4�v��V:�����|�K���3�=v�k�b��b��}�|���	�8r8:�9>&؛v�N�a:��a�h�P��t���1�&@zF~�+��{�PJ�����(���O�r�qC��Īo���X�+D1�-F����)l��eCئn���/��Ƴ�Xs,�9����c-~Fۂ�0�XM��	{���Xa�]bm�/�K�=h�c�
�@O��%���2��1���U�#&B?� �p>��=�Hb��0I�3K	�TbO�P���Q�`|�7܉��J��ܜ�8��{�z	|`��s	�ݖ���#�d��7>Ř|~����>��v�;��{�8�c�]���=v��>�؃��g��Ʈ8����#
�hh��6�D#L���6�4��c�&�1�*�(��cO:Lvld��x��f^ǄH�3"�|E��Rx��&H����tͣ�s�/n��t�*�cQ�DTE(���F�ھj�m���v�k��-vZ}����|l��v�X|��7X|��7ڭ�mn��7x|����7x|����8��΃�f� �R�����^�!�4�u`QL��2O���l�yh�'<��X�M����f��v��<ʹ	cf��6�T��nF�Q��4�o)���0"��&`^�0$a����oH-�q��ۦ�ZUcc��0cJ*
Z:��U�-%����E)]�_���34�	Bc�bv�ID)YYF&�Ta�Bk��7u�ڤyEh������~X�MT���{k9�س�C��bԦ�0�6��A~*��| ����s���S�M�aR_6|���C���Z���0�O�>�����0jSz_�R����c����w*��,g�Y7ķQ��Ї9;�4��C���\L��nВ��~��C?��eL��woВԒ�<�̇܇�1qSԮ�AKR�ֳ�d���`�I�1ƞw���`��Z��<������w-\��%������&.U��+��"�+b�"�+��"�+�"�+��"�+R�"�+��"�+2�"�+��"��:�z�a�}�a��}��a��}��a��}���t�p:l9�w%�%��
v�w�������;�d�/l�/�G��[,n˵wu�r�x��Y�.���m�$]r��߻M��|l�\���z3�mx���2�_�J����z��5�t��߱t:y��_��SA�j[󰜇j&����Շ���Γ�[��Px������˅?<[�=�׾��ج|h�;�|h\�yX���"����r�ֿ��a�A������|3_��x�)�2�g2�`�@6��/7,,5�(y#�V	
�����Z�އ��_߷��t2_�oܲ�2����z���H����{��~7��8g3�$o��ߜ��ov|δ�����7�l��� ݄��,b��o[��/ �ngd�����Oʩ�3��X��!%���M�+)
o�-׬��&�qFk@�e5���W��H��DllS#f���8)�,���	s&g���E���l�%~(�=���(�*�wx��{G�#�^������$%�uPcv�?|>:#dc�2B66D#d"!��Ѝ���llH�Tc�;��!�ذ�� 0��18�T9�!Y&f *f���%�֎��TU�ۀl��� نd#�Z���jZJ>mV�گ�_�*�������o~S�}=������	ee�]Y�W���±�[!�d"�G����~�X���6�?l�-���RV�2,���6<x'u�bɭjߍ���GY���fUp���=3a�����[��{?,�6'/�R1%�/�W�R僣Y^hҔ��:,�t������ŏ�O^cK�{;_�'�u��.L�G��\`L�ɚQZV�NW|������;�<�⍫$�pل�U�/W���֕�֏p�n�����T�֢��m)Cװ���+Yi�-�>H�k�_~�s��������P�9���W�l9��p��/�n�j�>��i�Ӓ����ۺ^���]٧)�
&��|�G�5��X���RN|���Y�2v��*fj[�t�BXMj'�rE�E�B�YX�U0+�X�˲�za"ԧh��j�5� t��BrZs_U5�]aҹʩJ��,�E y����K[/9X��Vm�|=y���7�~�p�_�}������͟�t���c��ޖ�D꛷~�7����ay�
�ɋ@��i�-��j5�睛/Gج��w_/�8e�����զ�L+��)�N���o�_�6��|�N��'��5���ok׬曛��C|'4$�%0;��I�OeX�Br�5�O-��4�.�t�0��)�񮨂�M�T�� K�d	S�� u\���Ckf�iɮ]��4��@��`#�ȃ	:�δ�R(�$`m�8ږ�����L�`:�T�"%'R�� EO�+�ʈ��/�}p����F�H���TJ�@%�N�cP��Le�2h��1�S�J�_[�jsڗ�Y'���"���u�Sn���W.�X_�^_�����r�͠7�:�,�iF�U1p!gLPi��|tʔ�3������P�f���U�'O"��>g����td~k"g�&��b=ʑ2�g�Q{�">�,�����M�g1KdX�<��s����ǁ��2�����eQ2��PQ�U-KY�u��m/O�K؊L���ݒ�+����p�+�a� �I���Φ�ə2lz)�jf����X)��*�L�b�H�]7�q�,˕ّE$VzF���SSpaiPaRٍ�i��@~b��(�5���m�H�Ô��r�,@�K��0{�|�5r�?:Ŧ�Ι���V�:h"�<*#뙫?�M��&h�n����o�Z(�6�[�����/����	�ܳy���wA�3����d���o�_�����f�����n�p��揓*���<��sMg��nE�I���}�������ۗ��w�ޤt�o��W����u�����i�-��i��o�����\�m�X%{�C5�,��]N�~,=�z���R7������(�C�QFs�[��)��#?�뛟��s��|Š`i0�Aײ�ɦE4��VoNS�xgm
S�d����i��7�P�qNp�i@kh��e��m�/p��N �a-����6~�t	d��n�;�>�0�1��b]8,y�V1�6���$�)zfYhо�œX}�@ W��&��L	U3)�%B��8�=��i�%k�U$f�O�X3#d��(���85ڶt�J�P0�y�`�8�D�X9a���~�tE��Y�L0��!6FƉ퐱�r�2A�w��ǭvt������`!�6h�N�>ݳ+��r��z��5T�����L�:�?�kK��H�&��R������L�{"3�Q���wLR�u~~���:?��iJ�:�(3a�S)���%��Xf��Oб�/h~~����-�4_�������3Z��dԆ+K9SS�t�l�6�Җ�'�����_�������~��_���MN͌+łsk1���Lɭa2�K�h�]�%Mο��������:;�mv*�f2��a��aj�)�zF�"�P����iVNȍ-��O(E\��r�
����m�;:�m�?<kӑ16<��7o#�6�Px�ַ��x'�4������w��V��r�[_��pL���o6�c�?�3~�4D��D��{"�	^Q�m����a�-w;/#�v�>�vAM�j�>��U���/�Ļ[̓�r��-���_���si?7/c�/�&��O_����fF!���\j,��4\_K�:lT�>���w���RƩ�|z=�pم����b<�Hf�� #�X{F�d0�(|�9M� �!cT�ΥsT�� ^T�B���	�PW . WHw%0lW�%��j�n��H��S�P���i|��s���Cό
���N��0��u� ����L�b@��D6�Q�-*$W���1�hO
�xd�3�=E ��&�����:ǩ�E��.'02.""30�.""0$�z� Fuܝp��:�jv�.vW W� ��]��t���v����}5QwG��uY�S�*��	����ژ`}q�t8X��FɎ��u��'a1�J,#�&U	����|����B�\�x�/B!�HO����$ƀ!�IP��K���+ܑ+D��ǹ#=` v���� QȜƀj����a-
�����ע�����"���U����Ť�/��6��?۠_!��z�+R��`� ��(���Q*ލ����{@�Z���A�k����������e0���c�# �i�Uh�.��,ȸB���!�\=�W�T�ɚ����������G�=m��G�^O�4C��.0��jٰ�� w��������7�۩�\��􈘅��C�q`���"�������9
�+��%��i��0QaG�OݱJ�TT�1��$�Pu������g���=	��Dh�	���Q�	�*�W��94^� I>���������G����"*�(0�|Ud�똀T����Pl-�j��|P�"�u�l�����V�r��s���z�J���Q1>���멶�}�0�}���
�f\vm<U"��^�t�*�<U�y�u1̸�����ȖK=j�Eo1L}5M���s\�xc2:��ڋ���GP4M#��Ga��E������᠘�?*6�d�26�/����Z*���ـ�t�g��=���ިb]����N��m��Q`��$'a�[�W3c��B:�6:����U�Ⱥ7�Ɏw��q�D`�6M�5hK��>B�����!�1��h�ǖ\Mֽ%7��Y§�ƒ�zC����gflh(6�������'J,ME7�%�^�w$�l@5���T�5��2�^kf��wL]!df� ��%B�Տ!����ِ*�2����m��}�7�9��}�x���%�kǁT):��0_,~n~t������ED�}���߾��-��ϫw?l�����Wo"��֫����{_��w��"&��PK   �D�Xf�� w ߀ /   images/04914e81-76ea-41b3-8036-a4ddbf8d15ca.png��ePO�-zp�A܂�`����-��5����n����� wN�����}xu�NU9����{��VϞ@)��(D( ��7QA9n�EF�(�tA�ㅥ��$E��iCLn�
}���0�k[��`0��������>���a�7D�&(���|���0]�x�����U����k��9�h�۴�x�n׻��x	i),���?�ºǬ��~`�b�10_c�	�]���ml�$o�T]�i3�TL��
�L{<_���y�����H��]X8�7�R+(��f/?��Mk�����)���;n�2>�ʲs��V`��u������o�`6��sI�o�@���U���Tgkn�lB?TI��(h/5�(4��^�+rƉ�'y��x��%��8�9.c|ߌ\�����d�k�E�=I7EW"���~hS?iB�
9��+)��(m�_,y�6Dɴ�r.E5���L,(BQ�ǥ�E�"���u��ǥ��;J02�q8R����'��޸܏�jT6��m���*)�0���!��u�U+Ч�l"yS���Ϛ��M��hHe�	T����@6/�U�4Q�f��';b'�3���o��+��˨��	X���a�Rs
�/�n���<��(�sH8��,��ӊY0e�[6�[��#]���l���"�+z7�䔙S�>�)���X{0������Ĺ񃶬ӱ�SK�h*����-9�o{^�45'���+�ٽ7�5�u!��c���M���˰�q�̯��kY��Mӏ|�%���������}�_1
C��+g��qZ����:�ee��iY�(��4������bd�y_�Dvw+�y��"�1��"�;j���qH)ٛL��E�]�!�Zp������v�c2�7�N*`�����0���]�l��O~�%�zč<NY��3a��x��&9;�S� w뽨��u�J��������p6؍�Q�ڋs_�,�7�(F�n����nMF��X|E ˿¨�W� C�:m�T�*O1�۶�����.?��:=\e$ט4Uc�me�7/��ƵG?�8m	blm����ӻz�c�W�)�v佽��q*�_F/`������V��7�^_x���D�m�F5�I�O��b��$�"5r�� n>�B�-䋓��ܧva�j$�8�����̩��z�uV�\�$+�m@�g�"�Gmw"��ο��D�u�WH���sV[z�Ic��Z��ȆL$����Q1rЪ�(�aS����AV,+Zfu�yu�ۮCĊ[ǽ�yR��p�]9P�� \+��`OS�*N2�q�ڼ]�sj�vT�W*d6�+&��1H*A2��-�[��G&Ƿ%��p�;���2�Fj�2O�/����l���t�٩A�?��Z��M�q`�
m�;�p��U�p��F��a"�L���Uso��C��������Wِ���-d�G.R����]�h,C�����Z�_���ث��͔��i��ѯot���1�r�������4�pG���J���/�����p�!��������V� T�j����uF�_.�/�6���ɞ���{Yl��bO6���]c=��	�ܢ���>���[�gb�u,�x�%foqċ�-S	9>iʴ`�.�Z������^(1�(�dF�$��+�0�W��#o��x�j�f��/z�ͬ�,�RM�?�$z�i�^�V�x/2{*�Wޘ�b_-�b»p�jJ��٨�D|:aG����๛3N�Y�7��
mi�b��CTs����?��^1}���%�E��ζf F���� &�v���Ƽ�)ڑ�M�� #O��F�Q�i	52,ois��9�;���2��6���>���F-j#�c��_���wu�EmyzfŅ�m��9[	}޲PB�}i�
~��ӄ(J�O��G����L�`�5���i~(�5�+c�I^�����%2��?{�+V�P�JI��d9u������_��������7�Yޥr"r�ǎlF[:z��b-��R>C�5Z��ŋ��9\ f|���*����FFg��+U�����+�nLA������X��*����:X~ng~��7]����Z ���p�W�AT��j{H	N�49 :�%���N߲?��n��-==v/�=F�	�;���7\v����7L}���c�I��jy"��s�X����-0����n��.�O��7�c�w����3��ԙ��2Y�`={Mb,zU��Tu�,HG�%�� �&n���C^� %)�έ�]�=4�Ty�+��_��e�DY�	��jJ��q�6ה@���m�9Ch}K~�`A �퓹��Y��L��ˮV��w�K�tN���顴��։��풬:�H���j�-�)G�%C늓���w�%�F�;"�-�O\��,HA�uN�c6D	_���ŻC�!��|�}�n�")�ʒ�ű1+M/i��ۥ)��>^o�~͖2O�)��}��K+r�pIx����{ll��%v[|�w��b�fbWw\���NE�A���o�A�ɭŚ�P�޲�_Oj%�A�M�k���ޮ��~ K+�?iv�f�!j��j�1��4�M�\�mov�vnoU�͋��N��z`�U��4@�Th�QF�;�G�h�24�E�:��գ��(����rv�ω�z���8[~,+e�s�៉	k����O�ݻc��h��/}�#M�q�1D�t�;9��-	�yYR�bR�:�~#��j߇�N�xy��ދR�J�TϿ��iD��H�c�Ar������|�[/<K$�	_GD>�r7Z^.�ipŤ98�~d��1���%�҉�*7��?�u�>1冡s ɦg�W��^�}�nO�����541{���L�����m���YB��m089c��u�A���Aژ?#F���D/e��L $֓�O�r�3, ����ɗ��^��wP�d��l�.��8�R��A��閻��q�][B0���p�ܸW�X&=k9&�:�7 ��k�[�[���e���C�M����ْt��VŪS���X?��-=o�m�����I�ĆgK�Жf��]�j���H�r�a��*N������8�xnY������㹮Bh��[c�gpԱ�f����ȹ�~�v���={�"���S���%1:9>��aʗ��y���	��:��$�rC:���U��T��+��?f`k�3�X|��b��5�7�/�c�4�Ǩg
��@�m��nŧ�j^
x�c7�!1��Ŧ�i/���"���@��{����H� �W�<�;yr��f�2��"�,�I���N;:)�����(���b`Jv��S���d������
wrX�`�Ucm�S�{%�� �J��I�����].+>���^���k�_��/zt��������ƺ{�g�b��ϑj��O��wîߘn7�|���e8�z��:�-�^D�����s{:WT�+6��ul����0���Tne�Ol�_�K�J5��Z�]�̨l���>o2"V���=�j��x�୶���)k�]Tu�q>�k쩕UGb}�������϶Y���j�L����7stq}�$��4�e݋<��;���������$(	$Z���ɗ��+�NV0m��uol����cQ[,B�ڔ4}%B��oN���6{�˻�!��RC��	�������@�b�-/��`Z�����O��.R#�ϛh]����3qy�а�{��Ľp���\�>��h��:W��@}��x�#9M0(5s�MEd�������1��5h������Qo|����i:�ʟ�e�S&6c���PB� �r^� �!�XM�Ds7��ogá�Z��gT��PЋݢꪋE�O:e)Gs
���f7�p��Ԃ�{��ږk����� >2��𣭍�X��<��Υ-s��vR{yK�t��&�����A���Q�
7B��#uZhՆ̰��Hzv������<��@��l���C��ј.���$�Y�a�8������ΐ�<�
��!��p��h�H�����f�<��v�UC��Z7��*��!����h�C٫N�U��w\��
^��
50X�4�������O���Όle���@�?v(=�G	>�[���ɵ)�\��S��(>S����|Џ����YQ�N7M�$F�w��(֧p��.��zm��C"cz_�n�eH�&
��5����m�1�����+�jTT����7���R�K^�"@�����>���
��Kt�z�[���9?
T]xbԵ/�^!�$�c67�G�M�;�-B�Q�Y�T�u�-�t��0��:/~�����":��fq��L�.�2.㘬s�w<�ш,�j[���@����d�:�0I��e����%΢���ʋ�O?9]���3Hg�UK3c4p0�UuηS-䲫=�bwa��Dh�9[y��`i��\*1R"��o�Gf�x������涱���J:&��6�mpx7�}(`�x�
$n���t1��p���W�agM�ue�Ǣ��lx_ױ�8� |�����Z�w^|z�('/t��zJ�P�EZ��ݤ՜�`�ON2��R�����l��F��X'�9~;�a��웦��4���6²\Mmv��Q]�Vԅ��q"�I��K/xP<���g�d�������[�X��׀5!&%õ��_���ʆS;.�q�楩4�� ���K�s:��e{mےnN�M��J�%��#���rm��ͧ���W7M����Rtf����-<o@s7@�"a���	p�3�Y�J��NS�ҁ	����N��(R�ݛ:7��3���-کmb}��,�Q1Er���u�!D��N^��2��C`�I��)��7�#dY�<"Q��*勉�1��(�*�q'���F~}��d�/���^4����?�7J{���%����R�I�5(�hF��iv�v���{��F��x*�t�/�g�1+�@rn>C�>֟�mV���l��R�b>���G�[}hX��y�ݶ�gy�(^ �tE����9�~}sbٲʆq��m�\�z���l���_�v�Wu�л�ޜ?�z.g��1�Gh+�p�ۧ�u!uwҊ\���]���IӉL���a�,�5�Ƀ3�d�yh*h�53�(�{nD�$����70���<�����Lo�ϋ$O��f��Ɲy�(�j�?:�u6�)�����Q}`���"m$��8�i,����q�3����vq�)7��w��\Y��޹�/����f��ؾ��_���/I��_��A�I۔$����V�i�^��j�L���g"(^(�f�k���p"�m��D���P���D��ˣ,p�,�f@p���(��l���β*��4�?i/5Ǐ�",/�!��V}�y(Mi Ā}��]&}�j���1O����M�2a��s��홋�,]��#�w��ʙ��bӻ� �~�m��B'9:}@X%�2}7	�TCH�x�����/��U�d�p��m{�|K�!xg1���3�u��e�#��œ$ɭ7&��){���'���d���]+�6�*����-��f�v,�s&8�1S����ݮ�dn3�g�Δ��&C	���YY�AOu�U��|��'Ռ�4�bѠ�˄�z+J�X!��˶s�V-���^��m&~u�zeg�AP�9+�Vm���׼ͱ(�Z��m��oU���|���J�|ʔ�cp��\�3?�2c�`8_����bH��Q�p^�܆qe]ي�O�\�J*(�MK���M�g7�;�����55&���G��7:��K�7��HfYW.�6�)X�%�e4�YvZ�V���}S��>���z��0DFNq�����{q�����FX0��R��ZZl/�m5Re�F�X���z�:ۅ&��;ö�o?���@�l�����6��_��h:���"��qA]/�Y��f�=NL��7���ݵ�q���1g�v�5köe
��5T�t�<߫�$Z�0P��W� b(r�~���r��]T��a�2۝ٴ���e�-?����$H�~Uey�6d:�"5�],!3�E��q��p�����oA����\����5D�5�)�_?yJ`��z�mS���������x����"����F��!L� ��w�3E l%�ңO�V�?��ݳ���H��D��3|tBw1SQ�%�؅,_����m�"���9+J�:.��mb� )QV�r k^n@X\rE�J)�W�����$B�<�j�G�D����u�������ZYu��_��X�X��Y?�~�.`i��abh��z��>��-_����#��#i��0�{����^B�}lN��ݎH�"CbZ翻��Z�*��Ϛ������v/�hK�R��Pk_��F���nN�EV3��S�[ۼ"���
���@kI�X�7�sw�?X�����zQ��񆢬�F�u�:�y�A�e�.�����8�EڕZsӃ��^�W�nQ�08���㔀�g)fܿr/l<a@1lE�6�#Jԃ7]�9�(�W�O27L{s����J�Vђ]Nz.���Vh�x��i�M.	/��9�{;�&�PM<�R�d':H-b����0���$��q72���R
��C�KjslxO��*�A=r$~,`Nle:ֵ_����y�d^_Nl�^��8�Ձn&�>�b�Ip��H��W���߄�Gp���∼{�CO��\q��I<�G۸��ׄ�E
	�Om�`��� �X�ލ���K����<��χ��}�g-V��ڋU��,��AA�D�����*!�}�B���G� �
,|rs���m.>�4Mɣ�y���17 ���l/�rp�����~P��g���(��X�:�.��o�|��[@���b
�ܨp#��EL�:
f(Y�>��:m��^�>�[�f�JP����O���¶��9p9O�?���������N�jY�b��xv�<�t��d�dUT_���ReԲ��:ߣ�w2�X����ɫ��P�-l��a�qj'�f\aս�}��f�y��o������<��K�=r]=�|amV�B�ˤ6� {���c;��ӒH�MLz�L@L�O5�S��~������~�06J�w��^C^bO�h|-nB#���È�MB�ly��D;���E�z6����G��5��Ċ���;��9����+��+=�,
r��y���Ϭ�A���J( gG�ZL��;Yb@q{��q��r�ũ��ғt�T3L�9��చ���̨�t�=�C��.�����
�/�BB�q}D�vsEp�^6/U��YL�Ѡ�;�K���eB�����[�$w5B�����n���m�`ߊ������hB�@�ȁ�O/���بuj";�.d�����RsjG��?�_~�A����d��k�r�4	L��I�* =����1H�+Y�c;U_�Q��$�i�ؤG��)�#���y��Mf;�,ԑš��q'�:�1 ^��rd\y���#����T�G�'I� ��t���&]K�{�x���(�䎸���օ_�ta���������੢V��,���K��1
�Ju�2W�ѼPÌ��z��Y�t���#�ghE����qZuW��8�I��u������8�&�3�$]��|IC�k��f&�K��[�KR�ْ�>U�]��YDP��Ԣ/һ�x����vZ�Sͨ9�hݭa[+ uPʓ�Ew0��:QD��0A���ȓ����T�/�����S����#�+�G�c\G�i��Yh��@2� �4U�g������r~+!��{҂�� ��1�Y
���J�4����z�k��x�l�X��Q��C���V+��5��QN3ܺ���YO9>�$�>M�^BY|�!��u ����okkW�gS��Z���?��:�
t���+�?��G�6T�cѢ/���f�g�Y�X���t�W�Kg�n=/��g��t����P�3������&�>6��,o>m,2=p2x!;�1o%$#=6�ܴY�[�z8�|�U��*!Yq㔐�;}����F�i���_����"SK����nSt�OT�\�-��yq:<��ă��O4�`�>�ӱ�� 4����͋� �\�w�t�94Gd�ܕ;?�v�������t�lj�N��5�hS>6�'葫=ܛx����2\�Ĩ�����ȩ�9�L�u������lk6��C�x]�L�HX�����*
�)cp��R�ڧ�,~�>/�����8��g^�R�|KB�&����͔�@�o�|�Cn��4�-����̊GMN[���Cܟ�Z߅L&�{�����Uؼ��y�4��Y���?��]���k����
��.�lw�7�������M�H5�Z�����+F�l@4�4=�6��:U;�E��/}���4��o�~ ���	�:��sI^Γ�-B	1�-uM{o��T���T���.�G���Zg�SV��j���.����RV�����^|���b 7�)!�9�{9��� n���/#�dRZT�ꭁ?&Af��\��7�����^@��f��E�1ŀ�:a�/�~�CHe�9�sy�]kj��zIJ �ִ�ɠr<yR�[�㖐+ �W�к$]��ݚ�Ñtol��	�fH�����e��ٴ|�dt���=['(Q�[v�D'U��ХΆ'�P���H��Z\Oc_�V��t&����`ֹ�}�TlbunW]6ú\v�����SW�֜G;SHb�)�K>��%�΍ބ��_�
��4�Q�����m�;��{���[}��3DYrڃ�[�������R��?���Ji�����D���U�_=� z���K�~���d�2�tj��e+�4$Д71!�픔X�l�c�/�e��5��|ǳ~��E�Q��ݗyS�e��K�5$���f���+�ⓣ�c In���UR��� vlP靥u��a��UU���u+�����f#mE�>�O�U��y�
F_1f�dnnc]�m[ZAߖ�< �%z����z8+�|��崗���/GS*��F��C�4,�[$�xV+x�
#AA=&�x��-�}��4�~Q�r�Ǫ�ifZHERH�ʍ,.�~��T]�p��iy����h����`	��p@nX�={��R�G9�fg8*���C���6���Gk�.꾪�f��x�A4a"o�v�E��TV�5l�_k^�xL"��<���W�MK6���/z��#ex���G_�uK����>=�����m��l�ᾜL�G��ZXFg��vx^���d�����-���0��]�N$b=��J�,����DX�:XD�*Y�:�ˆ���|�����^�2��*s���qڂ�Ԫ��܃��ȖY��|ːa#��d2�I:���z�);�܈U�p:"�(s0�!��@�1��1�vi��/La-�(�'�����{3����Ga���6��"_]���Ɲ�-��'�6���*4��6w0��!5j��[s��ڥ�#k��VdGB��K�B+���ՙX)1E=���e��������6@����E�`�yl��t�K��x�G��Ur��J����$µ�:���?�1	�65!�]�5�nmC�������>�J��|��k��۳�*(>������;����Z��lwTy��.��H��y�r�ut�C$0KO�z>��+�*�2c�����(&��wK���2���jBHd?mv�&5R(�hEO�,�{�J��*�<F
������%��!|��9���gny�8���[�VHnc�DC閈�5���臂1������	|�^)��\2��6���6g�V���@ٞ%4oZ �ȨS>��,�"r�X$�����M���х�^s�dh6S��|��)��y��+F�$�c)_Ւ�����jB�6s��^����kVjt�w�d��p��n�js���t(1�E�Ǡ�&�~ZA2� �2c�\�,��5��\-�q����y�4#�@i9:vN�� ���� a�T�G 98Ns$;�V�(�v@Q3�pb���K_�]��A�;';j�a����Ԓ�~~�W9Zwc�b�Zֳ����_��N��p�~{w+����u��(-W�G��'�3��
�U��:����ά��=V�_9� �>i/��O����s8��ͼ��9���6rV��O0�|���j���r�(��bG%*����xv�m��/�����b�w�b|����K��>��hF�wf�#�3)��J̉W�E�0�?h�SV��H\\�&���`���G�u�Q,�*;5�0� ���ɕu΄�)9�Qmz��;!i��c��-ڦ�9h���ZGn��f3�6�V���#b�]a[��4Z��`�fw���`+����^ �D1�!n}b�)�C�k�e�9�(Y^_����ߖb�����Uc�m���� ��Z�͕���x��<����G>�IsE"��E�&\>{�x���������)WZ��())�b�,�vՂkc��7��WP���\H����i���ԣ��'�T�J����9�r�V���u��$��y� J�\2=WL��>��m��an��jJ0g`�$�'f��\_i��6�V;gm�c2P4Y^٘Ț����n�Q@�3��\��b~Pg�Zn�P �{~�����To��il*_���~�dv�v�m�ֺ��h�1�zuխC�xݝ�D���Y�7�)t5�L�����VH@�K�gd`CCg�g#��D�� ƎU��1I�n���iF.�48z�@kו���c�`8a���5C�e�Fs���H��*����jZ&ۜ|6�*� 5�{�H���ɑ��q|`8'˨z�m=R����u������糶��]p��������?������	�lc(x�-�0`dy5�A��%��M�t#�ݜ2�<<|�hu(���z�?�F~������(�����j��L����R�@TS����,:�-So�
D:V��U�"��$b#Q����vd(�}�=�g�f�t�Vf�����?Gj�����;�.��@���M�#l�������B����u%��p�)��\!�3�H��Ӵ,D.ͺ)��@6+V�&���r(=
�(�|��5%Y7�ʞBƒؘ������g�Z1�S��,��sӂQR"z>�zg-#�z�F��;�L*�����-)?� h.�X�?@�%\ͪe
<9�A�K�Ԥ�dQ���uF��_M�g+����L��氶;�� �:g��1*=<xQ ^��}�v
����@��_�wMm�g�(��+h�n���L�8Q�B.�Q��B���\�̪X�c�� �1�{��vX��y����r�~��֙p��L��m���d�&
�]G�A����^���� �2��S���%����}���

��vd��_�8�����y��,����]2\�p&֮���O^�9�1�ru�!Z��K��˒�'��S�J����b���W��%�W��h����_
���H�^Z����L8��lK��w~q	��PV�6'��i�x�?;��T�p���yzO���@�D���`�m2S/Fg�G)��κ�E���QM]��^*Jt"�ToMbR~{��g�����6/�=À4�Y�<���驷��7�r9��-������A���3�F�߅�}���Q�~xH�6m��O�z-3�o�h/���V��T�:Xς9R�&'��
D�?ꈩ�Y`��6�xN&L[�\�mC�{��}��2�T)�{��gA��H���\��qs����9��I�&���r�8��J!�t�XF�M��x5Dߧ��ιLE*�RXzJ�Q^��$9�<��~Z�jqk�Oh�L>�MXhZd���'MOfܴBʝHlp*Q'��w��~d��W�J��h�?}�f��k`��3�J�1� -H���)�v��m����bYd�}Xp3���6��85��߳Wnܽ�-�Ͻ��O��{.�1oż�G9j�Q�/�����{�5^�������=�����{n��&�轰W��l��Y~��M��W؀��C�P�M�qqWR��J뉤PZ��uJ�(��BL0��ҧU<��$��$���-},�򼞮�O�����qه'?x��[� D��M�(�r��(`J���X鴛�h����CК��ڙ�dp�T�b�J�>EI��.,p��5?���T��ɉ�˦G��U�&��$:�8Eڕ�&��ؗ��#���-������ɸ� �=��|��@5G
�%P��"W������8I��")�Nu�k�u�i]����yY����_����wR2J}�B�^����F�4)Z�tU��_y�2���鍎���v@_���U���{B�~��M�Z����)���~�����u��?�=����i�/��{�_����+j���Z��?��h�����;�+R������E*��=��-�o����h]�d�Y��b\@|	�W�U�)��3�h�/��l�7�s�{K�{����P���㣙�ԇm]��c��9�QOӭ�(l��A^�M�v߳wt0q�4�[|l����YPO�v���>[���-)]�*J O�Kx���zpr2	M�XmmmkW�׏[Gp���E��M�_s��a��Z?��]2Q�q�o����I}=��	������Qx��kdXx͒���
ay�:�jQ8m��k�.X��֙�<��G����h�/�b�n����s��(��C�#Q�:i�����~���S+�O�R� C.�"���nc{�������M&��Ʀ��m$��!#eEc˫{�������Vf:��=���}E����%�9�Âq���d)�޿"�m��\2��0���Ɗ��ZYF�|�)�����s�"c�M]���b�!��ѱ���MF�V��e���s��'ঃQB|��ʙ�E�s�+M]�d`��޷��KMM�lj�	�?���9�v�������l���,Ϛ|ݬQn����B1_����s�>7��YC�����K��?��{s�b�/�7�?'''S����K��Ϙ4�5�QTDH7@�@>9= ��U���w�NtY���*Z� ���]���;�%�]�P ����O�ʞ�P��T�5?<�jD2�u� �a�f&lP�5�X���yx��SMu9�uj)
̌��L7ss2�C��/`$۟M�_mU~�.��\�QBp�5;�\[Z�e��� ��W������wttdiee<��S�tvf��?=M��T��:��� Ǜ����#o%|~��L�/<-�j�rB�5ǖ��s.��I]R�
���H�m_�|y;�*J��hWݹ���:۷����9y�}�*":*�[6��uk%< M�K&9Iw]:��ݧ�66��nZwvw����}.���:ϋl��,�ڝ��j�_o{�`A�"����%×/_V��~~ܱ�H�۴���k|���9������[<NF]M ���H8&�����乌�%�k"݀�'D�&}'w�Y1����p`6^%��R����p��� �����^�-B5�)'�.Ջ'��%� )I��|?&:z��/�n����������_���t{�%ɓ��	n��r�h��B�2����]��'�ƈuvw���D0��d4Vk����YZ�pq0���i����xI���flwSD�_-����iA�%�����9N1qAn�k�dA����^"H�Y̗3�js�Ξc��3͏�4��O��A����η��I<&.n}#O��ˮ����*��~|FFY<��ʧ�E���0#g!+2)�;���ȨA�d88>77 �%�|Ä��@:��1vww9��>V�~���^��l�*�? �4}y�T��u�pȦE����?�{O>D��4{�j����֌�������b�g����$#n!n��^��B�J���ju5+kk/բ؃���0f�!
ZZT!!�?�xP ����]������l��c�
��~�nfj�O(��uĩ���ՙ�g��S�Ϊ@?-Z-���|��($��@rn͍�ɓȚ�D����j��.n ����Jm�(�1�y#{lT@��
/9,�8�	�ϾLЃ�j
�ء=�&�d���!]��ru���c�줧���"HpÞ����i�3�(��K;�R�Q=������ 8~~^�|m�^_����I#D.D�;2������oM�u��f�����N��~���EheiRލ'C��c���s�m=��\X���.a��u����E=���,�M�E�5拖g����Ž��,T���ϸ@atH�wv�Y�C�t�Ղ�P����dY9c�7���&UI��T�K�Y�
e�b>(d��k/�@r
�T�����]=���ZG��Z�ء�&�����z�;��������QW�+x�bssĊ��K�윜�i-wV�db9���F����Q}1#�0���飯���e�n}����V��[��V6j�V��Toh��Q�� �g8����*�Y2|	;Ɛ]@��f�G� >Nډm�)�Y���t�m/}=��Zn�0�6��w픧Q�r�L�Ҁ9����InW_�k���˯�k����#Ԝ�[���`��7bۏ���=�=엑D1��lӈ�̏|�əJ��*+�����},T25vYc�7;;���`t1��r����8��P���!����V~w۝t)�5�F��NmZ���=+�m��7�-�qq��%ǝom�
-����y��ϘV"<(�#A�����k����N��� ɺ��e��~Z�:i�i`����Ø�F��B�1��=l��g��ˉ-����@��<�D�j
dX��s��Cx̕��`va��Ρ�D'�Y�0��ʙp������c�h������Ô�C�u����n�\j$4Ne5=d3bٽ �B�/��?i�	o\v�d�	�j�(͐X��1q�%��ϕʜN�bk���n��ige%� ���~�wx|&��nv���� �H���җXc�=sCX�,j���K�g�W���Ңa�W����k�h�2׉�ݜk�LQ���W�z�5�~�Jf������;�~�{�3��B>��t� �<u�����͝�E��J�ȸ�,��5�{+�d=�`@���3c?�n�H��UC�]#a&����ļ�~���L|GG�NIIICC�o$���|�5�Flٯja�1cn�H�{����U���Ѽ��8���3�^z\�|����8�~�N���{z|������Rpςq�`�.���/ O��ڶ��T�D�]����阜���E�y�m�K�Vur�D'�Ի�MR=Itì�3���-�o�~>`:����t𷎑)�p��d�>m�7v������d���nu�:��J����,Gc���L���+n[�dS0�6�s�!�"��q%��9���w}�yVܿ�V[�>�
	���u��:n�~��H����o�1|�!B�mv��m�@F`
�/'�{R^����{�Ŧ���p�b���yy�B��SW'	%�B��H:HO�V�(�u��5C�_��&����f���� �B��������y��wh]�;��۴a/���8r��%I�wt��x�1�1�Q��'�n���׏K�*(��U��2C�يz�C-�	{��jZg[��'&p���bVZ��7��jz��T�;CA&�%]]�|��^^^��c�8xx�vz�c5�L���Bf�Rs��NxL�޸�[�6��<�<"��h(��E���~sN�4=!nE��^cm#r����v��ĵ(�ğ�~m#FbԹcʔk��ʣ�}�X��e8�
3e�o�,�E��.�h !�\YMd��D懈�D�^KA/

�{!W�p �*�Q2�,c�s���MI����8���W����G�ŷ��H+����ۍ]Q�0���8�;dC&�a]+7�PQ�ҡ��*"�;���D�-��u���Z���k�胃���#������u���U���l3�{ֶ:��:Ԯ�����c777�|5e�;���:�*��0�䕨u�1�ؿHs#�7k�^��C�"�e����ա#�Wk����r,�Еm8���EH�Z|��L?�m@:+f�#u� �,
r��9�;~L��ݙ�5U�^��GNRV���S��.�|!k�#����aG=w�"���G��_�r/R4Ø?�@ߪ��i
jaVs�"�D��T� $]�+f6� �}a�z����F0���U��e8?��^d*��D!����-E-�֧J�t��Ѽ:\�O�R>�J�A�-,*�u��]YO����ET�������y�_χ�^/�<�����Z�d*����
��ί���H�i@���fɇ_z��ѷ�E]bˋT��jU,��%���O7����g�o���&��w)�����KQ�ؓ0	�P"��7T����<�i�\T�{��C�-cm7�&�c�kZ<w���Q�:���g-t'���,$�
L�nW#�-��\��mѢ�;:� �NU�4����J��Q�0��(�)E{������ֽ�lp�ӉsGEo�=�P!�ё`'� rq��]��Q�D��zF�iƞ�?UT��w���ZwR�e���A�m�U]A�����4t��鈒���˸�y���%��7 ��S��eϡ�`��j�Ե�z J'�}f<J
����D��2u��vU'���ϻvKx��-G��DSo������)�p�A�66_����{����kW)����&�������@kp�k��q:4ڜa������42(���Jk����F��"
 wK0�f��g:���">]F���)@r�k!U����� -�6�$Q�Mo��I���֧d�*�U�&��2��46��A��,��_d59'�+�W�~��H?z�>��bg����C ��ݿy�@_o��2�
���h���iRm6�*Q�g�� �px�ZI;t�H ��^=H�P��Lw(��Q({�p�LZ�z�=ng�c5�o|��*|��;���K�~��D�+�4b�-��a����r%D���z�&`��r�Ӷ?mM߾�QpdJN�����(�hDBi�.������f%�����F�k`@�n�F�{�ֳ��_g��/�����v^ɯ���-ҏg�.�b��xdhIBKJ^� Q7l���E(�ws�A	]�]U諐��;��_�~=�R�1E�Z�m��f�R!|�o����"k2L����\�q����v�	 "჋�+��#�j�W����:��:�t1�D� �ܑ�����e����g��&�in�z�"?4� ��knX_%R��s$w��#e�EbxY[/%+��k�{�MLnӷF����Q�Ϛ2�q|�Ƥ�3�J��R^��7NS�ޙ�3�0�wCoDʳ#���.����k����n��F�"*��	ׂ��HKS��3��U�V��XX,�u������������L�}@��N4H�y��VO "�#�z�b�
-ئ� ����y	��ĵ�,����!\˝�Nc3���;�'��������OS>b'��b�Z�X��cR����d����O9��y�3���U�dd��]��G�G&��ݗ�+�)�Q�O�����?M�Ί
��6�	\a4�gD��w�h��X�F3+?m�޽�x�oT�&��{|���_�2'�H;o���EQ�aԦ�R^� �] У�RR�c��|!��Io�;����U뺂��\�םJ"�+�����c�8�H���x2���U���<0��]^|b+a�,��Ŋ���c��x_��|�^�ӐN��1���".o�&<�؄�}�PέX6{���$��߲�}�^��g[�o��ZO����1���G����Tj�k�� +�Zv�W��?�?e �͒&����/��0i��T�<��P��y8?r� `�H�OCb�~�`��J��:�}~����u"#��r㲨�u��B����#!`t��D�5�WBd�~��4�<�ʤD�"�[�՟�ߎN������Q\+�K�N	?Z�����9�#�9�{��8@X�],w�.:+��E�7שd|҅�����X������ӱ�����/(L<]�q�"Or]���*x���NbNr$^Yh�/1��ۥ:�0���MÇM���b�"u$a׵%uf~���u��HC���ز�~�X��`��ja��b��# �kh������N��W�]�M���S��q�W�h ������ǉ���ߥ�׮,dXJ���b/�쵶 �>	�Ai���DW�U&�|p�^�-�o�^�7t����w���9�=�|�!!�g�z��~~i}�8�L;�=<�F�*�qoW/~%B��A�*�$a� �ДE�8/]����Ȩ"��B� (��6��`�̟[)�=g>Z��h�e(�E����!{��}af-�,p������7��pbF�M�ja~�ㅓK��Q 9�T`޳��Z�仙�#X���I�5/2��0���8��fdL��s3iW5��>jEI���Z��_-��Q�~dݔ}Ũ�.�A���8���N�Nj��t_�V�� �T��'�=��p������U���;L�4����4sN=Z�b���n��$�\���f��?��`���4� ;��޷����	Tl�|��eRR�$Ah��1��]�=����<m�)����)9ܗ��;�d�v �U���`�~�����r�I��9K]�sfF�}����g���w�B�w��4	��x�1�_��;Q3�o=n�OϪ�7����f�<�>��g��eK������,G�Y������^���X��>Dn�X���^J�s���d${��s���'�9	�^��Ƨ�$������k�7D�����[�1eT������ݴvla�nc4�?R�����ߒ[��f�qL���,5�Iǜ��C�2�S�Ή��N�������[��W��;�Z�����Ի����_�.)�ې���lo<c�3��7���oVڼ�-�ˍ����nĵ��gO�E�l��K����=��&�q�z�[e��_�����,P��]Z
�["��j��-������o�g�q�
e2�ߛ�+�)���F��ԜK\u(D'��]�DQ�_�M���e�f,�F��RhŹ�9y�3�)����KO���c��`,��n=@��?ڼ��؀9�
��@
 �>IqQ����ۉ�PՀWjꊽ��9k�>�͇Bz��8n�t#��ۘɻ$�k�S��ʠ���Nh����9q1�@�z�%j�ϽhW$z���soA�����)РK-�bM��݀�����N�q=��4n�.����"Zn���lŒG>Y8����8j�>É�@܉,`ᔢ�Uv�t&�z���>��P;���AK��ܡ����9�<$RW�����h�ܑ�d����SOIi�_ֈ���18�bmo|;��Ƿ� RyxȵO�d�+I�t�!J��E]zћ?�LzR �u�.4��(���Tෛ�d#�`�%�s���8��u���֗MUD��Մ�&�[Iv\�8���F�m�+"�Ɲ@�U�'9k��˞��D�&mH����bCc$gyV�Ρ��:�㶇w�4y�Ǚ�O�t����Ê�h��YFl`��'�#��!H;��.�����ں����9
�*�KN׸7"�ʲJ���� ����2UMZ�����rn<��0gII���X�d����񛽀'�H� .. ��	�홫،(��/�3sL��s"���)�z~$#C�a_�p1>�u��iʂ����f�!v��׳�1�J�{�%��a��(!�3E�ɒ���si�~�����j��pz8�/�z�K��r�#��Q,[�_?�A�<��5�Y�F����<im2����j�W��K�\P�G�r��X�NR�})W^Psv�_F\B8((�U���O��U��𲡂M ��������H�2k�_��������!'+9p����0�K���Lu^ݒ�$��!�~�TJ2� ��u���Z:��7i'�,�	��|n^sZL��9�|��:`�!J��4��f튂qW�g��VbOֿ�Q�i�j������?u�/<�81֐9�8��^mDZ_��v,�>_��t�4������A�ƒ�s�껶�E��[�^s8V���!�?����aټ;�t�Ur��o�MLL��=��Be��~&�bJ<�s}x���6K����
x��hČ�]��ܦ���Oġ˼�\���r�զ ����]W�D��u�м -Ze%C<���5��Q��
9Rz4[�)Ӭ��<���6_6�_��y<½93	�	fh��iq@�[=s:�	�%���ŅM7>��
��Ѳߞ�l>�/[���n��U�?��Ǻ�yZ��,���aV^=mu_��X�_.{R�S\�q���3���t��eʳ��;���9��uE>)����ϔS�yc��su<�4���2�QȈAS�+��&Xpax��7�F�ǂW��m���O�h1߽C����7�l��M~�����J��0{�A0H2`Z��W��z�e�Y�T�k��Jγt��g`re��s���!~���;�1X���a'��ĸ���ǧQ\��\�>�}�k�t��-%V��}ƶO������N�ʹ8����pT?�w������"����a�_�	� ܸO@��u�膨ʸ��~��ԧҤ��3�D�z�����bx�������:�2�/�_��=*4i�v��$��,�n��;�����&�y7��c6>��ļ��@���w$zF�my��K�|O;c��oz�T��|�"(�8:���q�7<sj�@�dV�\�V� :b�y2�pm���J��V���@j�}seq�yĶ�Z��WhѤ8g�n�7���Ɲ�$��X��;�留�ԣ�����<�FTE]=䇼�y�~�����p�٫M9�.�p*D��Z-��"#H�kp8���~U����CY��uw:�z�������G���o��ґW���&�H�Ӱ���q�y��U��p��kn��x�2k(��f����f��H�c����)�`.�����RD�sy2O�+.��0���k��kҭ�e��~m6�RtC�Q�7���Ւ��`�98�<-Ө5��s���U�cs���r��9t���fv΁$Ɛ���r���o	�^����Ȅ�����({�z�7�&��#�b�gA@����7���L��p����kk*��U��]�A[hWއ�P�� ��T�)Gq�k~�1��$�)7��f�;���0p�t%}PC�k�,���%�~������;XM���=�1�i(o�3*&	k�XrG�}�k�s�)�U�~L��)��.2$,666rj}kooo����i��,V�;q��Eӡ�%nA�K.�d�w̦߂0�i���{�r"л�5��6�9�����TIl��e����"�˝0+)����J�!EF`Ѫh�5���;��

�Zf��w$���h��,(���/��%��zÕ^���u���1��	88q�M��	&7��%r�~g��SA6n�^�
�7���oB_Ho�	�)�;"�o�����m"�t�FD�� el��!<n<�y=j7���qHK��nY�{<��g�s�/��85�>Y��J巻Α'3�|4����h��/^��KmRe��5e+��*iP[?U�^�+��. _6�s�ZQ01�O��c��&b}�Bcu�8� #N�ߍ�P��˸�fk�U��f����T���޼���� ��7��|�b��'���:Z�/�'Ab�D���7�ښ���
�!��:	��yV�����<d���Ю��0��I�c��5���F_����=��^>��1��`e;:�,��Zn&�Z�1���m냚v��(8]���䧺�f=�� ��Ҟ��.�R	j'ĩ��m~�Z�	��:�N���C�@m��B�y�~��������XoK��,��a���=[o����~�^)�O�kh���.x���켜bu�{T��(�~���R{:���u7Oi���m{��W�ڢ=���0��yi�L9�`��&96�YZ[��yq_[��eXz�2R���0��e���r�xν�	:���p����_2	Y@g�a�Տ�~�0Q�q^&��~DF���ٚ�$��O@Sg�G�o����i������X�J�'�n'���2Q�'��Н�ݘ���ǌ�7�C�
�t��A_dS��f����$J�ࠖ��S�3r���(u3���ef��0��ZPW���w�7x�lt�s|�R:Hw�y����ݘȳnmm�$�q�h���a��^�j8�vu�"ϊ������Ų6�ȓ��;Y�%�=iStǎ�U�s/>��g�[���5��4�;G7�G���?�<��(�6��.29��v�3(����_}�gnV���>�����]�\e�O��-��G�p��4��ͬaӐ��:gݙ�x�I���� �y��E%��ŵ\~��u���4�s��A&|������*�C7B�u,�y<����_�&S2ļ�a��^ ]�%,��'�v�L�� c�*=���:V읥�7���d�w�1��Y*�Jv���%>�-E�����d�8�Ӑyf�ϵ�/�6������I���S�MM$��$<���1��([����Қ;�=��U�IL���l�\_��~�8���ڌg�f�@y�R�>}�&|-^�A��;������I��Z���Y�.�<d��B2��e��xU&�1ߗߤ*0:�h�4\�$�$������R[M���⽷�����«>�~d�n���|�?˝�^h�7a�� �ƛԒ�ZKX��P����1��4I���J��i�)�S`a!2I@��YEe���I�W�����g�ˍ J��V?��5;�}2��KF�5����1=�y*:'��[�m��y��֐術�7t�}#���?�e��(��	��Ą����Ce�ky�W�2��c5��i��y\��%j4>�5������J,Ss������W'�kkC�V)#�jlv��X_�/=��y�-��d�ty��t���yk��u;��K�k1����PQ�Q��GDs5ḑz�*���x���K�x��ghK��:��^\ЏI�ۑ��cb��j]��>�C�]�vb8_��|Oh0�:��M����8��դOp$����Z$3q4���;�Zt���G�6@a+��v��/<&^
P,S�m��qt x�݇��ަH���F��Q�6��P��1g1	��/�x���R�v.vɘo����"�� �ĴZ����d4�S��M��ś?I��w��\�C�~�A�LD�)(��G҂�.n�i�o��d��)88�<]_�+�R&1�2�Eu��H|�����ɥ���c{,l�n�)-�2Y�l�9��99G�TG�����X�������X�5����0�16Ԉ3�izb��S�Ɣ��D�� h 	UE_?:===���>B^��R`M�[G���X�)Ľ��Y�~�2�("!�����92:�G���V̹�C^��u����\{�Q#��xQ�%�]V�� iR��<�vA2�bK
�N��p��lp�S����9�}E1FC'34 #E3��q�.l�9#?�զ�vϧ����c�	���d��Ac��,h����*jjH K�ލ�p&���Lۭ�����޸�U�ե��#�%��:!���#�:��>��6M5`o�qs��	�K��� t���,�WV���xxxhYX��[B��@�� �I,Xj���Cw魇@Qv 9�ю�}���|���uZi���4iI�hڠ�|�-,sg��43��-���� �%(���Ϯ������[���?����I4���u�]1Ʉ7�)�}ė�˺'o�W\�j��uȻ��-�c�O��++z��~BX����_\^�\�u����9�V�U��L{d���Qz�/��� ��l;��,�j�1kxy�.�c�������F�d�3[ZYI�����*�8���ox����r�ML~㰑����Q�w��9����"����p[?p��v��_D�3�q�!��`$�$k�P�K~N��w��\PB�~' �i��t���{������>��}� �w6r�y���o��)o� �4���&�Έ�������
����a�`�l�V%P�4[��Y�⚬�}����Fm���ދ�0[$ѮU�C|�������㠊�A�~�΁���Hx͛�����������
��tuw�ol���D��0>w��6�Lf�n3��,a��7�z���wKi/iit��T�)��[��v?
!�}�����G���s\�c,m���KF�.�-���$"��=�a�������𝈄!����rQf�%�� o�2�q���:�l���%b�hY�M�Hg .�l�(ߪ*�	�3練P,
�L��4#Qʏ��6�""0T54�����D���V>�ni���:R/]�}=rh��IJ��O��cKKK�u�����]��%����W.#I�'A��|4p
�Ǒ�B��p�A�	&O�痨��Q�1�ĝ�@��W���oz���������W�>����	å]��I4�,�IdC�x�pR������!F`u����g�T�O5ln�|�DGٝmF)��Y{���>Ǉ���r���*��U���\����)��/�?��D�w���I�7�9?;s6n�丯�=��6�#����^#*� $=S��e.�
-w�%T��m���Nw�{d/�����<�:q>ɃmPIʞ�rwB��˵J�G��@��"���$�<�~��*Ow����=\r���g���Z���k���=�v�ȱv��Y� 
�5r�$EU}��\�H������ H�i$
`L����A�a�H��nO�	ow��<:�t#oު�L�3G�Ȭzf���K�+�8;;q*<5��i���&ϐQ�o@�{�u9ib^ic����)��̂�n� �OQ���췬"��6޸r뾔8E�I�?����M:�ET��7���	�7�����--F��Pk�21��u�Np�Uc���(�r	�I�;M�U�_����i6J�GA��D�JQ�`��߻�m�l����u�-�9Uƺ��{��
���&�V���Њq�w��� �dE�j+~�'�<����D�%�;^0��Ũ�PLc<�Ԩ�ď3(�]K�n׹����E��>���	~����Z���|DF��=ſj��p�Z�y_ˍZ��$^O�?����wĽt�=��Fh~>�/�T�����~��%>,mLa�	A
�Y�}�j�{[��%� `$fls�ع�����������h�q�M����7��;����|{:(�5)3�1�$�ۺs�q��#�:����o|�N�����}��j�Fy눀��{|;N�M2dL9���(��;j�m��8��T�-�����Y��O��
�ǃ}�J�G䭆��.����U�:���[��R�J�A�yuMh��~V��%@-���ƀ�->���BL�xX�p4�30�
�FpF�����ˡ)!��\�@D�Ϥ�td.�$�ބ�]p��uT��{������ ��a���p�G�����կᕆJG"�J1��c<���n��s��ʆ�f��2�c�Q�]O_^P��P��3�k��h��oY�=p��Q}���#QzEq��91��!��-�-��w�ʈ�}IV���Lo
ͼ)p}E�5о~���O�ʹ��f�&�؆�2��#���y��7 "~�1����+��y� Z�J�#����E܉֟⹪|�׳����l���QE��d��b��xQ5_��h���>	��1�	��m��&01�ʫ
V�F��0�{�*�n>,p�)��A��GB"�r.5��lD@�?:�e�$�)֎7}e�W7.E�N��5;`�K�J�q��3M�F�,V��u����g�%��pth��~<����������u����v	]��"U�(��~�fFkrڣX���a��&w��'v�V֢�H�
 �%	W{}^��qJ���W[��?��
P0�YE��#wT�������N"�v��E:��l�{�?�r�l��m� �����@f4��5��a�t�,C�a��6<��`N��/I0PG>,�=�j�.��6���Vf8R���-���P�1�d�Ҡ|###*z�z�d�{ͣ�=��q�d))o�2���&�#�����}iύ]W�B�l���q øZ_n>$���c��훖ׂ����ԯ'�ҽ���Z�4V�I��Є�:�����ɎFj�����g�v9��Y����M��(�#��1��F͐��LD���}"�G���n#�A/>�њ���/��F�
��J�=��_Z��8c��::�[Sr=F�-w�іs�C�(�{�'j_��nS��̿���S�6��;��,:~��{ڪ��È�w��9�ޯ<rP��zp��2Q����8r�R����bn���L<��C���ȅE��8��t�&��'^��`��uI	�UB����8�>lϠwZF�A"K��w+����n�ج�����0��^6�&Ȫz�R;�^�t�̤���R��6��:_�����Ȯ�Y��K.I��`��/���ݭ���i�}���{o7���PU�<(=��A�'�t`�y���a�ivc��_��٫�C��2�吐��P�o�LPM��,շ����5����PMۉ�?nLvsc�3��b�ƫM�Aid��h.΁��������p��fְ����A��{���)j�c��~��$_�. ާ	ۧ	&qD���,����C�	<�����t��/R�:ZvkL�N�b��-[��Ņi	v#�!b��Qwᘀ��:���昫?�鞱�	�qt���_��L��tq9��3Y��Z��4" ��#��#�2>���~�ӟе��f��5�/S�J�#���(�G�;,o���#Ua�T��"�V�9�F��+�����g!���U�M����ui:����=�%U?�(�%����|PGT�R��E�PB�u7I0�Z<l� NLf��y���*�֏����v�a�?�&�ɝ0!{!"�ѩ�̶͘_��LY�ӢA����,Ӂ�h8����`ӆ�6�x~��.�?�����.��zL�^,,���]�ڛ3ڢ�VT�H%9k�
2��c��_���.2iP��eR��	��z̪����9dW�L���W�I矯B{0� ��{?�6Z�����F��m"2��%*��b�C4m����ۂ´��E�o^��V�`P��~4ى aY[d�����r1^9��������������[�d��.�	��Y6���Ft�ź���5]ٵ-��EwϚX��ޡ���1�/�F6�p0�*)�9��A��Q=�l�s�#N^��Nݡ7��F�J���թ�ɘF�ֽa��:���ZO%�~MMVqEE�ތ���ч�H��3'yy{''����7�[�@��Cn�v0Ը��#h�R3�D���+n��6=��������P�!���{�'��톤H7mx���]�p��wS!���ߟ+����5����n[��'j�T�9��E�TVB�����2	
N�L+�p�1w���ot�o��,1�`:].nF�`{����JY���F�m.G��ؑ�����!$�=���ZJ$%IϞ��j��  ��æ��֡����,Ch3u�rK^�lp��A��,��Z��= 5��U����DW�	�#��n��b+s=iN���V�i����)7 ���'Cc_??��'}J�����2�;POj�t��V*"�'��UHr���U�����������F�N���N�D�
wLM����9�����G��1���v���V�m��_i4�zBs:�ZC�fy.�V��D���D�1���� .�O\��6}���ϮQT����;��
�-/���K?b��6�Y����k��Ί #��C�n1zb���UUE�jχc�<�M���
�k��_*K�����$�L�-	q�U�G��U��93�T�o�#�i�к.��͐�,����1=M���ݽ�<&�Z����i�f���(�yS����Z�Z��n����0&�����SĶ�|$��Ⱥ�p��{|�������M� ������Yҁ�ˉ�5Z��
��Dq���M_�����C4�\�~!�9*�13yD��x�(���h��u�ޢ�H�6f�8q �A{�����r1����(���Q�OE~�dK/��c�Ͽ������jB��w�s=g��`��Y��=��$������ET� ��x�(l�ߩUD��.����s���NMM!4.c�@U4?�o� 	�ф/_�C�L��b���w��|����h� w������׫+%��?��f�J��;����Wh��/�n���#���^�&�;?��Ra�X�ZB�i� k�D�G�J�yx�E�&1[W̡(��$�hHa���X�)���^A���n[\5��>��ň�?ɬ�:�Nې�o�\a�p��b2�o�eQQ�G�[c'PDDD�T�L����}t�����\�a�F�f�^��)L$�L>�HR��°����j N���ОP�!N,#��EN2��8��;�P�*�HQ���޸�Jh�>.G��o"��F��������\��QԱ����.��=�PM�d�?$��Gm�f��Q� @=vW\�}
cE�X2�H�sl�y&�58�ꆚ����ۇ�O^y y9�J�΋0j�]�h�l�l����􏪁��J2���s��f#ɒ�/p�jjk��z�ꎞ(�pۉ���Lz��1�޴�-#�
3aʧ�����ꢍ�
Bȴ�N�O�7��8
uO�h��:���jT�m�����Cb<�4B�V�A�i͢�,�V�TFF^3��u��Ѻq�Wh���bK�Q�?q ����@�0x� ��T�VU�_Gv{E�ݓ��b<�č�bG�K#�(+�k�:�O��S��V?:4>>��>����>��kF���\�ؘ���bVtbI38B��{OY$iR�0xضo�G��3E������n0g"܈MF5׊�����JBDD���JJJrZ���p�PPgW�L��`��Ki!}�D��ؔQ�L���7;(�|��ߐ�����F�����d0��* �N���T+�x�n}Ot�I�DE�~e|�{1�拏��1.og��4�)��*�����A+I{���b�q	�pV��_�G[��ñ���坛��S��%)��wұ�}��):�p��v!�:S�t��V�
��D���s@��!���m:�q;�c���A���$�(���R����x8�/B.=���?���7�jN2%@�iA0�T�X�EC��#��)l+��"M��LM�vo?zE`��t���=�}��u��t=r�j�����	����\�Qʈ5^�1�T\^޿�)7�Y�_��X�&91Lu�ą����)x���y�yVez�"UA�$�)I�+���������_|���M�v+����2z`j�����>c
��V/��={S-*�@�	�uu�(y� E�1��3��qy���B���%�����ƙ��1L�d�c�yz��xq�0��C/�\���������:�@�N�Yw�߇�旽��Y�nxqm�:#Br��/��58+��P�EN��}|�+#|��$��sI�Tg��/�=Wpa�	XA�����ꔖ�P�Q?�-	��h�|�_���9���ʺw�ًnd��b<~z�d�$��Q:�Z�-�Ûg���yha�r�������Nv4D�r��B�gD��g�$1�WQ��i��, ҇�H�[�^5|4d�(�Dne%�9��9�.+�x��T���5���G"���) �@"���~���gҬy���+��׿�C�:3\w.�#i�`dwm�?��u#�/&�J]��<� Lf�'�[�����!��6r������`Ը�s q`���ƚo���2�����Q�_�OS l�T��Z�h?NYF��3�/�B�|U]_g�`��Y,.F�q&� ̂uR��;�vN1@1�u��q�	;߽�R&���L�,A��b�'D
m���C�.NN\>l��e�_^^V-�X�m�:�\p��/�yҵ�Ş�d�����Ǡo�`�j�,>-���đ�{�,X��C��K�eҲk:0D�@6(����%5C�# �D�;C���.�J�M�F�4���ì�[F{�F^�{���g�����A���R�Z�=�gz�<���z��1I�G�&	�I8���=��¶G�7��n~q@�}��
�z'g,���iܖ��}��+h�P`D~��-j������rv�7Pk���[��w__�>ޱ���8�x��ߘ;�Kb� ��*������k1!��{�C>�Y���\T�oX��	�܉�<�U�qC��.%�m3���|����zr��}+�<rV���r��țy�=�{I�$����c�5��XPwL��+C۩R�I��H#r�w<Yk�~���zD��2�b3Z<up!�S�A��%�d��g��b��,@����� �&n�ד�fil��3����JS�:��,�]��oj
�40/Y�	L�������l%7G��+a~�g
K��9��1�J��RU�}���FE]=q��GnCI>��o��Ux1m%>��62sy(i���of���'���䗑 %����o�H����u���Zt%.�~�L4�Թ
�Y��S��Q�M���1]�[]}�H���W���ӥ�-��OjCcc�l/5�Ը�u]��#^��?)_��Z�U6�<���4u���3G��L�:�9��4r�[���(9�}a������L}qn�r7q}z�-�-�Q�X�D�V;��ԥ��Z<��Sv�ͧv;����B�R.�هHE*��(���5�r�yy�Z�$��2Lj� �'�a�F�W����6ߎ���/4�f�?�%!I�~4��)$w+z�wh�p�c4R��,$Ɍ�ɚ�`dژ��Ѣo�I�`��+�^eqI�^'��ϛ��*�GY����e>{x�V0���G
 a`�\P��D���U���'0)�R�`p���e`��R5嗠�v>�WK*���(���KM�Y�u�|$ˣ����op�� ڏ�"瀂^	O�6��5��D:,F�~h0�EpG��c�_�'� �W��yuql������_�T*�'�<]��rQup�h3p�͇��즗ږ���P��|/��ImNw7b�I�^������\FH��{;5x��n	\�c�Ӂ�e��߹ �Y�!�k�_QWnu�~�����^�	���_���-����gg ��� 7#�ysssw߶����i�q'� �'���C�2!!���S\I���8A��8����;�at�%!>?��>�޴��Qǔ���C<,t9h#I1��]BVg2���H5��>��VUCo�Ѣ�p7�]��T���Tm��}��?ne|?,���.�����6�����az���l��-�xd�]��!�x�{�ج���EYZ<� C��nYC�~I���f�
��.�5j2����wt�YSN���|3�����U��v/�D2�$Bs�މ��y6};=8�<O�'"k7/t��fe��l9�+���	Q��Pa�K7P�t��VV���ӑjU�h� S������~���� �\"<!1WW
8� N�׍���
��nDS���J\8�W)Y� >�	! ;��1��=:�����'{�8%T7��G�?8�O)�L�U�?���v�CV]ϪG����ʎw���"&�Yض�&ss�B+7�{��u��n;f���l��)��3��3��&��z7���
Cf���?��K*�Ap��0y�uH�Z��Cz���̥J��h��H��EP�=���"���F�0`g���b��k��g�9ڹ_T���f^/��x�ޡ,FL����Ɍ�cL��E���&c�Ǚp�"����EQ���9f�B&X�ʮY!i0��'�]��4�
��#�~�c��4@���Fҫ��*�ֲ���^o��̔�H�m���Pwps�h�(�݌6G�,�V�&�"����V5e	b�㺀��O��]�^?�d����L��9w�;�����c� �K�"��h�_]� B	�D��"LT 8��^���hjy)��d��ɼa��t�#}�
+�]sE�4��h0��D� ��*4$�I:���,��\�����]���8^L9ј�	=2̥�y���Ѓ:O3/��AJ�@r��� ����d>h������,[�,ۓ�p����N�0X��E�
���.�����wa�`4
�Jn�)
� qR�_3+�" ��<.���N�"��&C��"�޽-�L������(7�g�lu7�����Ka��NA��TE>v� �:��Z�b�|�@\T �-�f���%L���������9L�e��GV'G�̦Qa�)b]�z��qd�}���c�w�(F��R��,�I�7��Y�i�qb�$�_4�y��Me쮇�O,%SX�;����5Q���X,�*(z��=���Lߞ�������l�Ksb����{<mi���.�����1��AQv73q&��$+�i��򥆞ކ�꾤�L�2QSe�4��&���UX�܉z�C3��(w:]����g9�V�mQA�x���h"aF�����
A/�#���ȥ�o��
x;���|�`'���)�e9�<�xR��)�d�U��93\cբ����oi�����vt��7�1�-V��9o�緈�+��WK�_}�=q�;�)�^�R۾u3\M�7TV9��l������:�Ǩ$3SX�bJ����7p�]�o�Х��胀������Mv +��Stu���%RV ����e:�Y���Xϝ5�e��$:$z�y��6���=���b���h��-�C��J��)^`��:OŒ��kۙ��G뺩����O��C,|�<�	���A��@3����K���L�=<T��ͥ�35\Xcߌ��B9Z���]�Χ^o=ݖ�z�H϶��5�x>�q��.��C_�$��VՐܳ����,$�������I�,�[EӃ�-�R$N��M�(�Y, �O?�L|�Hm��������������:ePܨ�{AT����:]��Úy�g�2Tߵ�Y����Y���<+_��B�����M�g@���U��� �z�j�,���&Ϋ�|���!��΁��a�˱��H9O�a��(��+�M�yhA���"S�)ߛ�m����� ^���ƭ{6�=�GR��=��8�V9��h#�Z����-"ړqs&vN�8������Z�\&{��R�d��N��` �E+ކg�+<�3`"�#^�ܰo��ψj*���r~�`�%�*ʉZ�|���bSW��EG�S8�w�,��߉�U�t������>M�}gY q��!�c���;?����P�;u Cً2���`Ե��ir4�LS����:M��aS����-�iY�����L�W��{������m�����V
c�I��S�Q��`ѵ�t�@t��{��7�w��@�d�;�y�I���.2�A'2

����Y�/u�EDώ"�<�0���]�j�Y���݅@��,���6o�,�����5r�m}&mҝm ��}���"�d����^u)R�H@����o��c��*N��м��!��0�y\�rv����Q��Am���0-���N���S܋Cqwwoq����ݭh��PRn��!�}�����e&&s��ٳ��k��P �!m9��J>?�<�÷;V��ێ��>����������1H�6���5�_�`��
bf[��Tؘ���D�]�����e11��U�B��5L�k���mX�������e>�Zɣ��e埩Hc����"iN��n2^�[xBo6�Q�R7�PM��aqW��K������ZWj�)cb�W!����P7���jNP���.y`�i:�B��А�����0��kQ��O�i��A]w'����p�{_��cL|͑���i�P����C���_&^�˥�_{�i�V�.\@���/ԯ2V�雿&V�Us�݆�r'��
N�eY'c���L/φ�ˣ���A鵞sR♽��I�.tr���^o�d���ѓ���>s<J�VNYM'���^�ʵ���?���!*<��Y�����zPn�G�V�3�d�ml����3rV�p	z���7�b&&�s<�Z◧ޗ��-['>�|7u�v�n���
��+��I�;�p�"{4lӍ����i�%��i���r� uK�إQ�����a^{1�C췆+a?��@0�#���$oX���PZG���&�D(�����Ks��n?	���f?>v��Ҳ���s�#�K$4���S�y��6��r��mWk+�e[0�BYR��W�$�Ȧ��թ��!�Y*�&��*��F�t�����Tuv����b��o����.A��ĵ~���6�3�5St%8�e���pj6a���`_lj�ٙ�S�f�`���T�7�ۿ�k��0�'�*���	7�mT�y~I��p�'`J�̾�e*+V(���4\�k���wc���]��ڬ��m G�`ͨ8%<�+6��ƣzB�>��N.� �TR�y�*}�����GA����,5ZA+@uNX��^s�_��z�]!�~�(���������PK����G����s^�F�f;��sN;��4�+��:y�4P�H�5J�R�"�=P���G�T��:H�O�;���)�S;��}�K�$樃���J�����ȃ�P����1�W/�ۤ���Q��@�mi)y朱�t�I�%�`&�����҈��Dܺ��v����拒z��j!��nmk�IGȑw%����6�A�E�DaB`Χ^�gL�7��1����k��K!���}T�|iH!.�Ɣ_��N����A�
� \�"Q,���Uq������`s�0��֨\�o ��LU�c��!�z�o���J��o�?��Kޅ���xb�GQ��Q$�<��J������/�i�V�r�{R9���Z��M����Ͱf%��1�D�n��_ɺN�1���o^�י�7

�}<GP���m��]]8b�=��h�\|�ug=r�����:����0� �}8X�a��L�ݝg�H���D�"�r�����&�d9M-׷����9y�h���s����ڇƖ�r�6~������������l���`��BU?���QQ�������i���ʋg����'�����Uf�u拣�@�����k��3���䩩���>�b�鯳��PN�`��� ��2 r�-@�an�yY�����
�ٸ|�~b� Z���K����`�*������ ��ęE����ώ�wF�ffL��.i�H>�b�4ڣ�Ѩ½Ο6��%1�>�ܽ@��:Z�����R	҅���B�"llb҆�+�� ?�Ü���F����5o!��s{9F1V�����Ct��ϕ�-e�nAJ��_�k���/0�6޵����}[GM�������3o��:*,�����������)"�60�pV9��{~�Ê�����Ƶ�o) t��`��-͓�K�Z��&e֏�znut4b����@G��%� �����Ɏ?�ܤl�j�jq~qN7<I�������u ����ې1N�Y��tpP1VW���ɷ���3P�0!ᫀ[Y��2;Cز2�(�z��Q������N�9A�_r��,�`xz�*/۹��0��?���̆c�=[���,=;	��')`ɯ����U7�����_#eZ�D�������Xt1A�Fp���\p����+��8�ά�8�
�Ҵ���>wT����
�^ޞ\��.&�Sx��I⁷[NAc	͢��wdK-!�+�Z�&�'l*���3Ų����M-��lbJ�,ڮ.M��QIh�Sq��_88՟eH�%�o2(Ra  �	ъ�e����j��⚚�1�e�*%%���%ǛГO҅��ť�++�L������b(����olA�2���-P)�_���d��,�!�����>���KL vG2%�;��ؚ�%�[��lbR���iӒeB� �w����p �����.�6=OiҦ~.ޔy;T��]�a�i�[���rf_F�P'L(�!���ۂBKS���^�~uy�1�@�a^w�M���(�	�g�7�	�YͲ�m�;JE��2�³��R���e�+`�WRN�	�}R��*QU����ވ�1eĢL��Ϝ�9��}�S�;���;��I�����l�#������>b�[g�88(����܌�*5�;+��,T����YU�{a��^�F�	�o�5	�c}Ul�9�&��N���i��@g�ϴ)J�#�����ce}�������l�K�|�㠯�'C��D6�څ�,8������
�L�Ʋ�A�|#���7�����G]�9��3]p�.j3�T�Cs����D�8���&߷��#/�#Q<P�h7�E/����c��">q�(\��t^� ���z5��pA1r�c�GL���?��i8�0e� ��]a�;Y���}3��D����x^�2�y`�u����c��Q��+�����0�q�U�V;%��o!��#򧫴����x��}��+^�rb��l��M�]��\�<�������OȆO"�*�j+-M��Ix'M��d�PO�F�R�\�Ō'3�� �9%���Je6����������Ѫ����VI��+*/����J-//Ot��ǭ����̥�o�z���ҳ�j��}��Ϯ�A�E�[G_}V���g~����	}����g� *I6"�T�"4Y*9��=�ߞ̙��Q�) 3���;W�KOT1M��\����\0`�Dx��lI��oA5��@\���>���@���Q9/�a�ٓ	T��X�K,ę�8j�;nDBvr�-v�Z�֤;u��ہ� _t��/�R�xXʩ��L�·P��eIoq���X9&��x���(a?������^���Y--|]�'n�6���<昧fo�E��]�;��2���+>�~�R$�T��i۴�r5MM)��f{yu�oC6�Z��y�̴d��o3us��q��"���/x[�	SÊ�e��<���$�a1�2c8w�'�M���Ք18���Ց�ϮIЫMj��ZX�3���m�ñ�p6J��`�8�/�����?z���-��d-���������,�3:w,omo��ʪ�������D%LB,��65�3�P�Yו���ّZ���F��q�A&	r�����]�C�/�aI��Yr��� +e�x���g�tb��n� "M�e[{紘�W����u�D����|	��}�W&P�c�a͑}+�����;�w��V�A�;�х��>����@w�K��\��&�OOKJ��e���Z4����)�wl�j��,-��m��h������»w� ��q>�A��S@C;��`�d"�(7��:<���ޤ
�	11� �i���rmν���"�o=]�5{���w�t�h5����(�[xF����@���U��*X�rG�D��f$��w������I7�JO���:�m����f} j�Q�N'��Q��B�xͮZ�JV1�ؠt�8}-�����ܼy���>ؾ�8�
p<Jn��X����@ϊx��W�lx�#�~��R��FK7�.y��pw���qnu�'QNfh]D"��RR��M�ӪȆ�F��'�b0yn^�M�rQS��3��/��i���؄j���j�'v��{]	.㿳�U�����6���f*�3e��J R1��]$|�p�l:����|�?�=.�E&�*R�-�W��r1���΍�<�|A"��7��/�/Y0\Ǉ܂���"���[͐н�X�V�p nˎ��d��@&c��Z���y�uす>��{�,޽�ܾ���+��iX��cXR�����S�Ն��j��Õ�,�
�DA�n����<_�� +]��Zbnp��\.@��Oe������(Sg�g�(�c���,"�LNKk� �A>-�}�ϗCz�?rz��z�fx���wX�ǃm�;tT�D����s9-����޻�O�������䤵�C.��9���'��H~l�zٗ��
+�V���S�޽D�gEE�������J�K�����5Q:ڮ����ox��,���e��sS9�,Њ�������������Ev�>����+w�&P�햇�Ϻ�`a�f��.��s\N��ƾ	Y���|��.�o������4����绮��u�󨛴�o9�:>�������/��A�:6�&%�3&@��9.nj�h狶�$�wGd	g��p�c�J�m�����_sb+�\�`������J\[��ֱ�@�mW~aم���ZA��*�W�CK1�D���:���"�Z�D�zI�K �W@AE��l�P�<�A��H�w���ۯ�x;���e&:�H&9&]5A���3�4��s�C�N�PZ��"w�L�������Sy�����~7��������G�8*"Ѵ�6A�<2�X>�������Edn���ѹ���4��3�
qW�B>��$��@x��}�{{,�&�	#W/������̭��[���R�:Ŷ	`ኾ�E�l�?�� #�P`L���`�5J�B�s�\��b'�݄K{8���`�T^E�r5�����!d2SS�8�&�������v�v:\���w�f������֨ús�D��-84 >�hY|@LoXϿ}1�t��PҶ|J��n`�0Ί��Z��7����99���_`<m���@,E���Q������ǯ�	D���'��A��f�ts�֥m�[�M��[=--D�=�=b7RGg�3�8a!ҙ}����F���~QVn��L�R7Q�4��yn�W���ҽz�<�3=��8x��%�A��А���p�I.���گWp���]��m�̲���ի�&I'ǁ����T�/=�ؔ�PAw6_��࣌A���=�|Ls��H.��?$�j��ZC{ڲy־�u��j��V�%��N�N)ΔH�v�='y�:YAJcu��܋U9ܖګ�+��	��8�gk�����so�\i���h�E�s���W�][�>��sO�
�x ��<���v�}��t���F7\f-lu�JU�vn�6	�b.��M!m1�N���Pͼ��cQe4�LEX�q.Yf|� ���������n�e�H<�h��Ih�}b��� �`��1���g��J����[u�����-�.�� �Vo����cmo�b��B:"���w3y�'Wk��F~�nAwPN�$�\�"��b�Y�����&���_���e&����η�2�s�ML>���r��8m����
��#_w��o��'�o>����l��E��[�$�Ҍ:���Tȥ�&g9L������"��!~tW�Y�ծ8r���G_ˋ��R�["�[,�J��!^A����.�D���]SJ��\���y�J�J,�8#[��r&Z*Eq��~|�/�E~�һ� �b���c �T�~����B~��{Ωn���}�tD�!��6%ҡ���>T`��kg��y���?\h�XZ�/�� f�R�SL����URRz�A{����c��^Q�tq���f�-p^�3��D G�F���>?߼N���8<I�lW^acm�=/Wb�F���۶�Q��P�W�|f��<�F?"���s�=����UB��RD��,t;Jߝ,C���_�Ҩ�;.ġ��YU�+k�B��zjeE�n3��Z���Ն�z��n��u8x�ը���ݧy�z-g�w�)v��ᦫ�2J��H{�v�jv?��/��/�`�:���]�	9�3��I����y�Ma�K����ld��.�S�o-��V� �Dj u����<�{F�t6UN�9�	�9jR��)R$"���$��|�R�9I�S>�t�:z=Z�@���Z��m��G_d���D}�@@�KS;y�k������ �F�K�Y�����6�Oqχ?n����:��|b�GG�--�y�266�/�>�L�
+��+g~^���
��r},�uk�t�*oh]�p���K��荄i�����x�q(Y������� \V�%����HWW�ɠ>�}�YY�}��Cƅ�x.�&�+���UX`3��\�ۣ��D"�$7�����_�]̠�DxA��_�	A�����g`G����Ck�;� ����<]��^5�+ix�z�a
�-M��k����?kjrvD�F���-@�̐R-�L9�?��)G%>쪀1.�	���紐�ѭ�y��z^2AQY�� �������<�\h����v�C��	}&��s,�Q�R�� Λqn���)�0C�̈́/%��͡��v��svl~6^a�Sf���]�E+zj͑��x7�����R�$�/��;�� /\� }����x\��A>�s����ZR[GO���e55���R�3o!�e�j�ŋ{F������i�3o���L�,������^j:].c�C�*��S���:\�n�N����^${,+�fJ�C�0�;�TV�������Jħ���
��7�p�]�K�AY�u��#?��<M2h|���5߱���|���C��.et�g�&h������E6}��mWU�ĥIW���������x��"�����8^�x��71R_Y� !���P'2ϋo:�����9�l��A:��� 
�!Ԝ���cXO�̭EH����U-H�f�SEf�cYƦR;JF� �8�ل�J�l��l���QU
�7�>wf�;$kQ�\
xd���|�.�/��t�߬-�*�tj�{�K���}_�
�*�,���	97#���)'���,'���,
7f�oyF^d�b�S�_}���m��V���!��Zga3�_YX������U��±s��4������'��j3Jr�HE��� ʹh!סZ�^�'y�=����#K�Ty|:�2�:��-娤�$���"~i���,\v�_^^^PU���W���e 4�B	[��#}tY8��vL� O���9h!xi���Ō�����CX+(����@,�O�:�~�E{E�c�:ґV�Ng�ӟ���:K�Ih�p*�\�QՄ�;'c۶ވ�-F͚h{m��qs��g0��vr���0i�p���A������A@-��� ͬ+�}OD�vծ���?a�I�Xbc�i9J��Y�O���@�mK�5�Y�~ �[��f���[�����|Cf������d8R��ӟ����X�����n���Ц�gCVOT�Ml3wd�nb��De�����4@�ޑuZ�Q�P\�PǓ=,�6@gm��65���g���	�>HNMu�����/@�(`nE�SxB�j�>}����\�4|��T	��0ͫ� `Al����Og[��Z��?�c9؍�Y9W����ⵅ�d>�~�e"��wK'���h��YN��|Iϒ+�Q7l�>��y�GA<h ��t��!�ތ���G����)9��YC_��(0iL◣��g:*/���<���Rx̬��)�Y�6���-z���bz�n��2�t��y�0>p�V�$�BD�G���o��[���r��Y�dz��;�[�~vy>�8�W��?*��d�J�j��1_�����}����-g?��d���]6c&��=�(�1P��f�ϟ?��@�?ut�eN�.�p����(���z��\��,Q� ����(``r�!��)��(�b�����3���V��{�l����@MY�x�����Q|-^��za�#�9\��4��/�����l����K��>����܏�q���i�Q
�*���.����~����f�y�8F  �V��X��3��_]�,SI��@`�	= ��p{�/(�lb���D<0p�(�M�%ͮ�l�-p7-Zi@�p͙-��km��p'��\������J��>C��D�)b�|ݡ�I]_�m��m|�u��n�࠰�52^�K#�� �@pgr�ǐ��G��kJ�ځ7�n�s�B20N���	~��vi� V�;&�g5rAĻ�!
��p+�j������J��堌%��&"J�^��~�K�ءI�w2P��6!��a�����>%�:�QV�աU��
��i�����I퍻�dޣ�ĺ^�i�B�����J2T=	�7�ÿ��E�کFdU_������ ��[�9��@�#fBg������V���s��_�<�{��RQ�+,ԑ��e� b��	�G���u�[�o/t!��;���|~U��f���!-����9`��Nfqa�` �1H���+m�ֲ����y�SeY�3.V�PƵ:Wƞ�؜���X�*|�O�(�^�2�A�]�D�@��6��e�}��V9-��^$�߻�|�va��s�7��~n!�۩i��ٔ��������]�e�xe�zo"'_�jP�Ÿ1���	�=�u�Ntirb��Q����c�����]����3-.Z�R�
�[1GY��P�ѯ��l#  47�h~��+�R�H��(��X~�j�'zԱ���G�����4hz�����Y6aϰ��k3��-���?b�c[��͡3iry��0n���w����(H�Q����i{b�A�9J�͝ ��5N��0�oy �l,3_jT�h���o��<7��ي;^Ts���2D�qы���	���'z�X��>k\�RPl(�n���^�j��=:�����^�:���� GX�Ͳ&��[Qء��9N�����ڎx���͏�o?�k��������u-q'�G�o��:G�x
\��)��,�hy����o�]mP?8�g�rh��WP��uI�ϊMz&n�$F���{��D���%e8���Q:-�K/y�g�����s��A�κ/j&i��ѣ�N]=�w����Y�>ޫvKINq�(�s���o��}(N�c^�����%hf����^�#��(���c�r�{��o�L�W�'�)]����<%'p��`cn��	.>�#�\YY�'9t��Z!;t*f�'8���@�����>�s
�!d�5�����78�$zs#U�:<���ț{�ڮ:���j��V������dAR�wf������M}�̝C���`�Z����S��)ԉ1�)��"?�砊G�m�<�g��q�8r�]�����>[��?�zv�KZw5�@ü���ԍ |�B�Ӟ����Z�g0�H
��M�y�q�����,Md�Ω�����`:V��6�>׮"���`^$��	�պ|G����N�{��l?��r,T�C�ɯ�h�ԏzb���͉��|qR2&��20��ͲK�@5��;���_�z6K�/ڣ��)6ǂq�Q�Y���Ӓ�*O��ǵ+�x�x[���:�p��N]:�s�� ��z�/���jbH#}j�hV���������H�lLrv��঍�{t{]���u��k�7/(xr��g�ɲ��w�M�xh�w�h?��ph� ���ê��Y��F�J��}�1��v0��GʛV���ɯ�R�y�?���#���Ǌ�(�� �N[̌5V5]�n�a�˥*c��r�nWj"-W,�z�c��CǞ+w�Nu��@ov�QD�Q������|�C�˅;%!:�y&K�I��>�RݧÓ��� q���,��*�fFX` \ٟ��f�h��Va%�ï z1��;.�P��A�+�l;�/���%�1o��>8����1�e
4�qS��'��z����%�.������U���۫c�S�jL�6����$�Y�� �<7&�F$o����)��Y�O�F�_��<��Z���}��{-�������Fe���o.�ouϚ�/.�Z����>�Ʀ�N��{z!n�e�t�ѽ�8ڌ�v��js�{�����<�0���x��w��w�������>�'�?��lk��z=J؋�Ė&n�4�C'a�bK%+X�i{b�N���'�R��݅�>�;�����<v�Z.�	A���۵!�/�+�(�)�A /�{xd�=�?0y*���$�GJ`�(V��1��0�-�T�D��]�Ĭ��ɫ�G�I�\�Έ�%gڼ�3�첊 �辗6i_�;��u�|Ki���3۝74�^����U�oz+	��d���캦�=�}Nf��ꊷc��֦!ûD����m�=mZh`Z��"����9�0zu'��N��9<BAAk
=����{e����|G��*�[O���F����/�����v"��v�9�mTݜN�9�����2%����3�!u��>JC?"8'<�=����۔�y��Y�Zၰ<��j6�W�� �S�V����ӹJ�<Ծmsi�KުV�Ӳy�O���I��-)ht�:��h��>�Q�b�[(�ָQ��� W.��	U@��_D@��/!d���v����{ =>n�����F>�گ�k;�X�?|�̣}�8���������?@.s��h3�V7���|i���0s7�j��U<�T�,��1Cm8(_�g"��_�޸\�4�z56�<��?��7h#�~�<�r���cY�����pT^��f7M~����h���n������hi��k��\#�@��baļ���P�Ӣ�9����z��I߬����:��b�0C�g�~@}8o;�V����:�D�:�`j6�<��^�G�bl2���|m���$)��q�*�K�O����3	�u=�>qEɢ-v)`1P�;�M����P��b%�W�����X-r�T���%�&	�C01�Ju�Ԙ�x6^����$43>_1�&S.��k��`d)r���'/˭�1��5S�Ogt�pP�Vn�u����𴞊�|�C׭y��oRX(螟�35��"-�ۍ�.����f�2�Ҍ��4V&>�U�
�H�]�t��0e�*������Ѳp�:��E�r O�Sǘb��1�E�
���z���r���Duf��7�3�W�Q���K��~64�\{H�X0\*�#>꿡�^
!���R����,d�$�`:��ip���L�tݮ*Q�@��a�ln^�W��:{1k\jG0��=�����j'T�\�2�����{��>,��8�G=Ic)���-V5l�����1�B��'��E�y�Ap�$�x�t�8��Ӵ���O����p�j��#���^��9�����tiQ^1�-*8^��!��<�ϱ]�LS<|"<I,���ne�]������m5ϓ6[.�>{y�vW[�U� ��̬�ӎ/ʐ��Ԙ�����%Oh��(GTE�"� �
-,ߧV'q`�(C�(�����Le�!�vj�����bX7�A����+��7� ���:!���mxu����]�*���f09�S�Tݯ@x�=b�8ǎ4�4Ƈ��t�u@�L���p6:�֌�Ǝ]��9��
s�<OB�(�PUW��l p��mUM�x�,j�6���j���V�"���jw�������,�fmU:w�Ϟ\�~��F6n
v!n�R���I��V~Qt��B���٭�X�Z.\P���� =���GX�*��NR��KW#�}�+�8��9.������0T�˗Q����<�<G�|��v���>䷴�[eW�����Z��3GQ�������'U�!jU�-]9D]���
EB�>�Ӭ^���_�� Z#*�T�T���֭�W;3b�T�{`���hw���cw�1�M��yFF�0ƚ����R�o.�W����ww,d	�����Z<�Ժ���׼C�?r��aBqt�O>��%�XJu!&��VO�ri�mjz�}�R�R��5a�����(�";8V��XP��U�[�����gP�<�M�h���Po�L�-;20��l��I��jQ@�ȼ '���U��˽D[��JA�۩Mm����%&�I���!��Ӳ#��=K8+�0��8���j�<+8�;	�:ʎL��Q�ϑ������E�P���Ywy��8�B�W�#����6g�ʝ���Y얖-�*�ȍ�6+^�gU�;��-$5u}>PBBb7#lx`��e�f���`�VM4K3�b�@]�G��,���2)��n�š���-���б-;����-�O���_��Kh���P�9a]K=.��ݏ��߬C�D�?��L�x�h��N*7CUWee���F�(�A�}W��k��Ɓ�|a W&���K7��ޞ��Z ����H�y�Z�~g8|�T�Q���7Ρ��aw���+̰�w�ݐ�tUa�aaBH"�,G�+���O9N����[6.	.��2�
����U�z�6gT�R�Mk���@+S!��(����{�V̠3I!�QO�p�Ƚ�ѕ�������z~�%<�rnA�������fy�q�^�$//<&"�&~�����4$a|c��9��A������0Y�w3ոV��g��/Af.EwN��ߥ��\!x�b�`��ꪆ�XÁ��H|�1��E��dg"�y�^,hdw���Il��qz&:�O~�ܑ�ob�A�#��Bؕ��bҭ����D
|OX�h��$#v(L"��:�|�>��R*�������=�1n����YSC^&��8��ut�A�y7l���A�il��P��,��-9��V��H�+_T��fm��Y�Ll�ƫL�0i
����7�]�����I���?2n�pIyEz9B\6��n�Ӟ�{�s[�$Wu���0^��̮�G@=�z�fK���u�NvŮS
}�Ҭ%W�q*��Q��o�ƪE�Bp�����w ,��C}�b��CǨ(X�*��*��jP��J%�\�I�84s)m�d9)g��]V�K�l���3��v��>!XY�@@g�@+7o���U33J6���2B�^����<�����j�g4��V��������;7=��&AU<���-�U9b���8��_�񢗼r���$=Lx�6��"y�������u�<*��p��{���L��7�8*�%		�ik��I�*3��1�$Fl���'Gv�^�چ���[�H�1�n����}�M�/�%�M��L�vcP��7=7��=Ӣ��Y�c�-���B?�7��Y@y���&&�/��|�����(q�
��ޑ�`e�L!�qϴ���D e����'oJ��W���_��JX2^�x����j���TN?�����Oh)Z��9�!�δ�.A����y�%2y|�d��CG25[��N���~��ȿ�I�Ε�6��-.��3f;����ߺt\�����	;r��h��չ��z���"���� ������<�������>?�=���۲��� �Bt\�M:Y���k�'˫���:d$ȭ�(�w}HhS�ٹ��=5j���(4T��(��GO���b:LFyӆ{��%�<H�5T��-��d�W.�b����C%��[ ��G#�X��ӄ� ؔ6��CMbu���?,�U�|DX�O����bkvDW��3@��轌\p��n�L���9?���e�P;��,9��W���nf����􏗺			[��U���A�����I튊�����}�����.�����[�Y������u&���cJ�x6>�a ����9�G��\)2��®� ���M%%��M>5�H���|x�����J|;r�0���OaPQ�dF��v�&j/�Hp�S�?�@oII�!��/Z�}W����:��6Gkċ���"UKc��,m������x�'��XjMQp22Z���˛���s�����v����^^�ll/�����gyt��bE��܏r�/z��o^��kAVp�H��>>�2u�fiX6��a���x���j"\�4;��H�ʬ'--~t���oSӥ��I~�m�����9��X�M`����J{��;ٓ<O�濣�&G=�.EƗƅ�X%�,M?�
D�-fdh/ �;�@,xS8-�p�Q̎� ���w��Y�&F��,a�%6�$\ �I��,����N�;���&%����&@U
��J�ș�+.�pCnjm������P����<x��Җ�f�(MG��>�u�G\B"ġ�k�X������5��^ ����7��f6�F2NuZ�������&u)K7+9i��U'��V5��_ټ�8�ӌ#iI�0b�[Q̶Q&��Ԗ�d��A��d�H�dե�D�������3�����d|�S�W3�#�xG��Ue�e���l�*��#�
߶�`�z�|g�9�Ux̠n���'�١��̦h�A#�D��O���ʗ�^=�:;�p+qwc�_���נF.R��2��D���-�����ż =M����i\\�].��L��K�!}��������y�K�2S��`�
7Y{���U��D��݇j��N�S ���F$d�ho�^�'�MM��TF���:@9>`��	v�GIx�0�+�]�
k�^��,mv�:��ݪϲqƧ�������)�b"����xٓ\J/m{������*;MH�E�>�j�����#��w�J9��5<@sr=�,C�7�2',-)4��Fk����J�ݝ�?�6�0c!GcBd���� ���s���@u���S-48t�,�`H�=a�ϼԋm|�Ce�-ý9��`������lz�5]���������N���Y���M�??<�������Q�q9En��f����Z$\][�ٝ]�T�{|\�ё%�����߮g����>�B� \\���ߛ[�o^˝��dۋf�k�W�h1+�jm��BEO��Y��ac�؎d���A��ꘜ���}� ��Q�ȁM+�F��)\���u���[�����R|d��OI:|�Q������}�Ƌ�/J�/x`��H��~+�>@Vx��َ���:\Ѡ�uwe��iTQ����
��B��'SܩL��w���������_lt�&���s�o��1���*E��VjU�=����B���ȏ�fļI�sðO?�^4{��lk)''���mom�����iL��O���w��MI����c>���b��W��~tx�1��@��/{<vJ�1Y6�[�0o���(=�X���w�z7��g2}��<�X�2��z_W�I62̐J���!��y	��ThXh���G�L�m�J��5q[ J�`ee�Ŕ���ͫV�ߟ$�]FG�uj�cm�8�G\�E������,GaT�/ҙ��������B�	B'aF�~Z(�&3���P���j�HR���S�{6n��|��6S�}K���z��,p*���D:��+��=-�}D%��/C�L�u�}�g�XP+��t�|���z�r_'�z�.�<���a���s�ueM��PJq�eL�!{���J�$���W<�'���#�dQRb/��slF՛c?+uX����P�<�Ί2�h�a�f��%I���]Qzt{��ӺLO&(������'�=~��Tx-xBYx����d4��q����i�*�7�D��><�"B�po;��tn#���['&��QCI����>�,a��gJ�N�)��Q�������V�?��Q��=1Jh�^TI�1��\����`�ɗMϗ}�p�r�L�SP3PI�"i��mrP>��χ�iCV)a@�̡I ��=��U���#WK����B�i1�i&�@�Cp^�XP���DZW;I�p����M��+���NM-�J��+T;5��U�n��'2J��A��sA�ɢނ�*N�C���?�g�o��:]�e�J2��O���IV�-/H����Ux��il������W�{;�9[��j�R�hF��g�C�H)6��81#�>��2@�D�' N"q� ��VƗ[)�C;1����0'�4��o1m���)/�h������z_����}�gz��C�؅em�'a�����1���7�����<3��Z���꛱�\�%;m�F���v�RG����i���kv�R�q~���ڢ��a`2!�eb�� G�����i*�^��+�%K�lJ��v��i���R����J�S�)|~/Oj�%��-��%�U}7X������  ���Z��C1���	��ft2���{*���[���r0���I� n���J�ID1�ί/B�Պ�@C=��C�L��L,�{7�j"G��k\����	Ɍw6�R��,W	���*D��>DW���i?��N3�����$�&����@�8��]���\pc1yO�d�����cE��e>?���ٍ��Z�'��3�.i�vS-��#�g2��2�(��v���u���æޮg�/�0������l��p��y���b!��x��u�g$,�\��O������GJ���*UMm�4]T���V�h��A!��餻��t�f%%$FHwwwH7#�Kr��������9;g��lw���<�}����V�;��1�$］��.���gF$\������mb202'�ŌHywt�+y���mI�⾨Aכ#C�ͮ���ضo!��k��oxʆ�{_N��[��5ix����������k� �;E	04��{�I���1g򞎂�>�)�@�=F_�7��|�jZ�F
�n�\�������P}b˗J����ZΏ�ر������}�
ԟ�3��Y��z@�;.�zD�:���=$�0��_�{���3s�
^�i��|�[�K:!F��ww�,�,}!�X���E����#}��\L7�� dh�K˟�`��T�����{����+�k����>��ݸ�-_[$�ΎAǃ!�V�����B�X�?�f�4����Q(˷����C̮��Dy��i��F��S�݊L����B��\&��d+�6�o�x��E>�s9M���^�:�G��/�6�$}��8R� .��	�w��qYUQɧ&*o} �����J�@���$6y<�`��. w�O_�T��q"�G�Oh���'3�V������^��,u�����J_vF}u�y�.�*M�5"�K��8���K���}��b�<O�x�y��%w����%�lT�d����Q�OE�2��\7�A����u�w/�P���F������v��Ӧ�㊉����'��;)N�,��]*��4��0�"��P��\Dz:ں
g:ڧ�H�[Tg疆%	Ъr�h�J�4�3�_����OvXOvh^q�g'��c��k|`��.Ѱ.�^}ҡ˳2֣���'{� 躰hst��Vxs�R��s�p�o��}������m�z�s��.���YĨ%b�T�<�/���u^k%��D��[ԋ�݋��
P�.�|��BN�3��� �wp�[T���d`DQBCNhF��:�^*�S��r��e��,=tPE�a��[��>g�3<����?k �3k�vlluVN��m�P���,���O�x�]��jD?>l
��ʨ�O���l�|J������F�x�<g�/|��q����Ih�
~��XV'ip��!%0����-��^/���
a�SSc1ٞGZ��o:�g���Vn8+^��e��>��K*_Ź�%Md�~պ~�	��×��@�:z_�R�3��m
���Ǚ9�c~�����[F�9�:/]����͝0���m�,L��U͵RK7ц����!?�1�P��}�ȣ}/�'L�1��Z����TU�4xt�Ȍ�(���G&��Ϯ���lѽۏ{ݝ�N���Jvv�!��h{}�%�3�N�MN~�޵�M=�8�Cȟ*mN�89�J�8���`F"��B�Lq��C���̪3�X�����%v��V�,�:�sw��}�x�̛���j��+4klz:"s��POԢ4 �s�����hz��`�v��u��	�I�l��+��/Ђ�}�#Z��=S��	�	�:��ʷqo����ǐ��6���{Bf��&j�뢎u_eq3�4�D�&��B���(abK���5UU��Q����>Ef�����+aCd�m���Ӏ)}H�x3�l������W\�vG6��6�Ϸ���|v��
�1_[	���r���ƙ��$ xoI��Q��M�[ı$�e3`P*��C%���2��T	�m��ϫ�����3�{L�sOt�	N�&�v�ra9HM�@{\��a�)���_���'kmmݾ�U����_�X?�T���P�k�~��y���+�� �0�lC��)&,ׂ�=��K�gj�Yg½�.�¨k���e��=O���w4��@�~�,�w~�n��@��FP& �&<gM3����kUO�-���uæ7(�:��&P�J��]ޛ�>��1S�$\|{��*Zy�:o���'^�$�#A=&��2�X.�����0_>��~z�>T
����| ��֠����زִ���>�;���Z	&���BMi�}��l�1�%|zrjj$$&_�H�����cBo��pkkL[< 8k�k�K���/�#�64y�����g����T�^���"�w�A�wW�T�'ԡ���?�=��5ш�M�����F��
���D9zП=�#����}���|֗ �0���/���h��M�\�9�:GA���2�U�g�
l?"|u���n	6j����;45101�� �1���%�M8�|}dhhH�������V��uŊ�{W���ۋ��J9�7ȹ���_��1��jqU����7�C4W����f@�?n�nn��x���G�l{�8"��.\F9H�|���X�C��f�����|�?!}����T���������yqa$'�P3�z
ZU�����T���iY���đ�}tJ/"ˇ%�g!�ᣏ��w{n�Y���?����ǡ���=�j�ķ�6��կ�Tm���Se>���*�J���M/�B�Ӻv͹�Q0��
���>���B>�&�5��P����(��z�����h}S%�Xʡ^3��22���8�)������ػ��X'�I��1GF
�3`�۶�E;n�T}P�Rwg$z����n�E�/i�}�r�Y}I�M�v�[vw�/���?�Mčb���eu1�\NU.���Ǿ��Y<�P��=�B�B��p�?hC�w�'d"�����CT������wh�]]���A��K��]A����1UUU9]���&�*�����qL�^�`�s�� �v�OR��o���t�]��ixW\�槮�چ꥓�S�������̠���@�j�=��/����p��汅��k��C��&�l�^Y��L���MVN���Y�ӌ��&��g��7e-�/��-�Vu����F�r|˂�lɸˌ��V�O�i$C7eu���hf�T���=�R�cdĖ�P��[��q�]Kxp$y�۵e�@]�-	������-V������X��)�T��|����RQU� ��R����t��*oՔ�W���ջ�B�
!���4|�#�����+�It1!<��N��\8x��Ւ��5�*J�iEzpp0{����(p����'�vO(�}~��w%|s��<e���l�����%�}��:����'�NI�������2�#��n��՞�4�>M�
��h��J����#�.��O�A
�w�F�A���j�}�r���t�?x§�=�r =ٷ7Ѕ
c���F�4�W/���UϥpC���x����1� 9�ͪ[�F�
�"�K���5�&��fƛ��Ѧ�7tA�e�_���]�wV�ǷA�>�W������(��
$ܥ|\��W�8.;jZ�F�@�@�̰����A������c�7��+�_����j�o�����2Yț,1��#��-��釬�H���ק15��y�7;��z�V�g#�&=�i�֤H7�6Zg�?4������Tsn���d��F����%��3\��k]�zu=�Ю��G�]�@��\��s���}�n�95SH4�ޢ� Us����]"K����lEڤ��˧O�e�`�}N�a'�^?��f!�PUW�RT����4�^n�YZғ��~��-o<{5iwH����������|���ߠ�\�IR>�]}y����;H ���ո���*��Tx�Z�� �-�X[��'��E�k���.$(��Wf�'��u�ghQ(�Ԫ0=}p�~}�+�z�`kB����;�My�N�f���яp���J��:�ac�>�Z]�v(˳g���j��/}�������l?�(2kkkء6�������/\~�pݏ����Ҿ��
u���6���	B������E�y?|1#fh� N=��#]w�ʯ�s��Ռ��Q�a_������N%)�����; �����mN�QݮSS#O�5�=��ʳ?.U^;�R�ӥ���_�&�c(�z��C�N��4ꆭ~��k��ϞH����3�U�#���s}��-Y�j!�U�12nJ�f�T�~x�_/���D�ّ����Q��l�t�f��&j��!�/�u�9U�����?���oi�^B����n�z�m��ٻ2�'8�y��;��Sm�9;3?���jC��ʫ�j2O��9o���d>T'&[��B��֎����Wz��73뢺�+I��5n��������S;n����4����vnB�wwN�=����9א��+�̦"���$a����\����fq�;g���y�x-�����S*�u1���<��q[�=��J�-#������F�UX���>���<w��]�r�j�a�U��?¦��Ѩ�8���� ���X1�.^6�4�;��t��%[��$��s,��M�tv!�YU��X��1'�u�N�2�m~r)%ܴ�[oZ��Ւ_
��z,k@w�� ���i_5,n_�]pi�?� U��u�_|���)�<f���	Ȓ�;�>�3���(@S��\�deS�ɀSr�^�i�@�g��r%{����ք�3���ȩ~��|F�d\�Jہ��u&�2������\w������J8��^���9֖�����p֮�,l�T� �
K8�a�zD@�7o1!���2�������}W�P���λ�A?g>w4�n����rr�^$�V��
QnJ��֦dм���s�J6r��Ŋج�m-�̉M�h��%�v[��
VWcqW�Z������1�|Z�1��V!�\��i�a��b���/����Z��3.��?Ώ����l�O��N����� �ׁ�^܋�U� g��.�4=�/�>o.�?�'�w�bS�h��V�����L��a���$04����Qe�~M��ތl�n
v��Z/=_�F⯧����L���}o̙7N{llI��B�1�,p����*��h�M���=1���L�j��j{n�F���(�����ޱ���{��tǡ�۞>CC�6��r��j�Ѝ�=t��"�
��:�!M�F��SŢ�1�b�y{�"^�<k����L>���@$�}�J��yCxf-��j��r8Y��2�M�=^�w)ի��>M���,**���x��~~���iٶ��}[���}�T�=�O	�=������<ĳ~P�Z!��9�D�+Jh-ƽ����*^�ڶ��Ƭ���a'jO_�i94���>VPC2�����q 앬���F7A]p̧қ#�!r�,�pG�l�&%i��Hk �����ٞ��О(,�(`�#�J�U��v�|%�\p���qS�#�[V�K�8�N�(�ngH�	f?�-љ��7�@��11u��OZ䔔����AD�4��<��&c��;�at1�k���|X�� Ga�hW�ݫ�\�%�.�&�=Q�[X�uܼ_��I�7&h�ݏG�
R�;h ���X��.ЬV�p�S�z*�.������V0r$��7Y�b�g�p�1[�LS�d���řC����<fbԎ��jN%�<uQ�=q1�0�<S���~ăTUU9��3;x�Ġ�1������φ���b�/\�<��'���H�h�$w��U�<u1ޅ����os7�!��{$8���ؑ���e>�iJ��T�Â7�%�!OP�W�$xᅖ��u�L�|��MfQ�W��\H�i�[8ƹ�L���mm�ҭ;���b\���g����&�Z��Q``��� bڲjm�dww�e��FiAN��f��%W:"UD'�=��|�t���轥�?�6��;^�������)G7&�Q" �>�eU9��rF"���QrE���(�;�����I��J�߉�RÁ��8����a������̓�aV}��!9��Bx^-�i��Ɩ:B�t�e�|\If�g��[�h}�rw��`������:*/�?�:�L7/''����D�M��ԒP��K�W�5��\w$6935U�s}�����d��X���m�2������I�P��{)0U���
q�;�M�ܒr���2�Q�~�ń8A��6&�m18�"�u:1tWo��:&/�=F��Y7�B���7��i�\��F//�g�i^;N�����%>�\`d���K���hb}���
��30��LBB;	В#[��4����1����vt�2���pI��'0��k�q=��UJ��d!�wr�X����&� !�����+-?�/�Х�`���1�M���K�I�S��$��+^���'3��h�������l�RH- �k�,N��C�l�݁΍k�]Ë��7��G�fJ���#���95�0),�^n�m*�n��R66zJ������k�\��
����X[7<�c/D�u��d���6��R'�0����W�
|K�o�E�)�@dHf�SӁ�s��X^�K2#~�Ĭ�]��i�ÙR��C�b[^@�dੴ���%�'�@)\:����L�@ї�����&��޴g''��Fm5$t=x��{O���Ɂ^)��/�?86����p����jk��I�l^A���0����R�Z;g��\��<i�� ��E���'��'�"ѓ'�&����ţ
Ip����19�7oTy�@k��d�Z���@�D!>�[����3ϟ�B�k.��+,"r�%��y��Bw6���#s�y}�- ������H��];��A1�O.-�V(j�X}rD���
g+��Xv]ftD�mgG*]� DB�����U��d������yƭ�LF�A��v�%�1yє�ƱO�{�5G��,�D�,:�!,�a�v��N���+��n&������Ha�_S���.fl&I�`�Jdۊ(�����bmƐ�U��Kʡ%�q�]m�o*����<�(�`!�����=y9��̻�\π <H�t#=1����W!}ĸḀ����5��Rd:f�ٱ�sY���<�	z9X��r�n4g�
���o�]'r�	i�O!�\fM��vQr ��������l���e�N�li�������doGLma.)����;��5��Q���طzϟve�܇=@Ȥ-r�G�����G/JR9��pςp	��]�4>�����7ѯ�9���J�V9?偔��ߙRH��֐�Ā�Yv���[A@�����qe�c"i�������q]���?�~���W�P��(i�to�e71��A�f�^�ˮ嗇Ϧ3�����UH�n��DXGԿy*�NZ���pᾥ��T���]�)0}��jX��{�A)�1+�;�Ų��V�D����3�����eMC�h������4;��S�Q� ��ڰ�^|��������f���i;�u�e��{�fA�WXo��8�4��%ZZ<c�W�����iXs�eI���R�2Tvۿ �ur�V\&I>����ȩ.M6%���F�ݞI���m�ġY��];�"�X��'W��G��O�:�V�vy��f����a��6VI������oV!*�a����!g?v6�J�	�׋?�9+d�L��q`�x��l��Sg�X���)�f�%��  ��|��'q��hJ����B�?4��Y���}dELR`Ȉ�\E7���x����^��[!�����#��ȶ�[��k����y���QQ��Kjd�������oYg�_�	T���K,�7%=�$NF�[��<į@g[
 ����E��PY<r���w�U�O�Z�|�sw	\Jr��5H�9"z��x<�-���^��m�!��ٱ�/�q۸Ysy�:�ڎ�_�w�뫼~;0un{�{�x9,�Ȟ��[�pt�s@�����D�M�*G��;cg��59h�-��Q�8q����"�A��q/��<�\tQ)�	"�̱N�ov�C�-t�nN���%�^k�'tk`Z�j�Yt���f��tp�)Pɨ������Zu񻌽*�/:5���;M�'i~�t��{�\Юj��E�f�����	i2�%��1����TI�A�*��?-�s�a�*@f���J����֐LG
ʱ��F�*��R�1�^`{N�jT�h� � ��F� v5~9[۫)LbT��;2Uq��DKFor����Qf�n��o��wn̏���c���X@�PO��i���?VU -�1�����~����R�������v��>��K�, �,a2���MJK>�̨�3+� �[n3*)�{��P�<����c�t��|�����=2�
�R?z�)AE�d��0b�`\�ȝ��gk�>c���I�3�6�0�J)��f��.�/EK)�ό�����ND� ?�C��n�)�^0���FB�͒Y9G����p2<�-�����?��/�����Xo!c#����g4okT[�ULI��(�+H�9��|��3���^ʬ!�T+9W�I�ݜ�\3��h	E��[��IAYZ�z2����e�['V^"�L�jz��C.�_�xx�[�4k��"�2^,q����J�R����gd�_����/�
���O'�!
$/�����qe�IÞ4_��:(����ڇ�Rϥ|��k��zK���#���9�b	�ˢ�����fn).f��@��S2�,���hu���yjO�ͫ'�J�+��mK�� ���t���l������	j+�1�ň�G�ċ� ��D2`�+�:�|�u�Αa��9̚T��U�F��<���
HlgJ�S�żwk��Њv�]N��
	�fCՒuT)�I�#"���7P������F�O5��؄� ��R��H�=�z���g1bƩ��'h��LD���ɕp�������\I5�HM���h~��R����������ݦ����r�K��8 �E���i6�4M����'|�m�P�������>�����;&w@@�(��>)�e�S]!!��ո��%��̘�90>?/��ec��
�9z8�w����`�!�W��U�<���R��ɷka��Yq��_���"����X�� �ۂ��$W�i�	�6�圆R�Bls�o�I�U^���S�`�&�7�dϿV2&�}B�(���W,�ߴ]����-�:�"#�c떇��,��a�}�p�r�q0,;����'��+�狩vO���R�����҆��Ll��?���E�u�����t{�-�aN�Jׁ?���"��N�9�Ƌ�|�)�����v;�*�tg�
�35��`0ŦLgE1|��1��A�<)���SyN�G����C��V�&���㢃�i�-���1z3�6mʖ6�_*_^�;I�>�aem�}u�Ǜn��9�I%�V���,�C24lllqI3��h����r�Gb(�p�-���H��=I���i������w3˝��p��M�Q��ӫ�Wލ�oV��l��z�.e��!10S�)��c��Dd�m��)�h�N�O���M�ؙH
������Q
L({���J�%D;
�C�[zX����O�A{�6���2j?��;٬Ӧ�X���?�"h�����_�m��ӊ��_33�ZZAf�������~���2L�=f�i$MuTi�9��mvu���-�o�:��W*�I�o�p1���[����.�.��+bcb�����M���ǯb{m�'+Уi��<�����!��]�uaU��`�� ? "�x�X�� ���v�x��}���S�]�O:����
L�Q��x�"�ᆺ�f�wr� �lv���ؖY�߳HXh�3�������=�q��7)/.[22�v���4��0[>�X�]����]�YN���J�R�^����W����W�گ�9'�C�X��:����YcV%-S:�V�������j�|R	%��tl\�A�cw)kRny���}�#%�(�6VV�|��=�F��p�y��Wpoˋ��D��e�q
��O)�V�V's�F�i���XWc�K�/��,`��^+ܝ�bX2���K���]���#�lʓ������@�dF�s�Zp{�\2��L[鉴.��S��	Vu1��@��r�F����n: Խ��s���;��X?�JM�D!޳��			a������f6",������\��������S���0@Y�nQ�2��H^�~��w}y�}�~k�A��'K=�<�z?�ϯ���ޘ�՟�[>� ]~�oR55oC�����mq^�j�����v�v���x���l��E�iSVf8ζ��y8R�z��tn�����bi/�>�9�i3>:Nf�"��8p{��l!�E��4j�8bK�'�E�.��Hw+��Xc�K�u6I"�Xӯ(V��L ���|U���f��.�J��:+�?d��ѻW8�	`V�O8��Q��ZS��xxѓ�p�-�F�G�
�~O���e�� ���oȢ:C^�I�"D{5��"��Ʌ��> �N�	��!M���z|�3�� 4{1�N+«1&�3�j�țIoۯ�+C�_c=�(�p�'�J6�=��}����#�'���Ώ��������\,3�� �ˮ���A�ٌޘ�ti�o��{�����>�p$���7fë�l���
����Gٹ�~H�����-��w��R�V��6Ǻ����~Π��4@f��^�}*��RIO��{���� �I�Ǹ���M����_=
��7������ߝO�UO�"���Z��J˥(ֿB�X��7#�6 F��y��xu6I� <�TXo|b$$����]�m���"KV�o��	1����yv*c�֍u|�̱���|kdS[�m���(O?���Q�x�n���\�B�tjK��++5פ���OD[�#g�o�'�iR��I0�&�a�}fqVw��A�s�x֑!�X�z���L�	}�\/�q��'�7�� U�t��f�]��%���G�	��'���))䂂����SE�E';Y{���Tt��E��viV%݄vg^?�p�/LH
˯�\�`��bЧ�t{:C�#N��)�ߤ�c�i	;��I#�s
�k�;G��$ ٘���w4�����������9PF�³Om�G���V��pm��(u�b����߻%e��e�8o.���0�:��,[�O�E�.������$mZ�
3�r��K�kSK/�����M�ߚDW�����������;�p
�GImG�l`��o$��Y��6�J����#�;����~�א�����wN� c#'�H��ѡ:c�d+[[�x��bD[e�v��x�ܱ�ZHekvLZ��}���̯�MU,Zp|Դk*�ۥƝ�ۑ���g�p���hmަ\���]��hG��b�h�z��;������~g�އ;� �X�2FVl��ֶ �{��)�49΃MT��E�Q��d:L��H97(RQW����<��t�u�?��������l{F�x��Wi�nt��T�t`0�?�z
}�4��m���G�"�
a����ƽ��D]�nkj��@Y��1��=��+�M��Э4ةl�en���G������md}����T��|�c1Z����2�7 �1,�:��?Q/�7�ݲ0NOO��$\]]'��_���C.�EDDy�Y[ë�zq�`�Y�s^�˧���A�m� �;��Q PrƤ�JZU�ukk�GkL�������JM+�X7m�t	�-�����M���:_*ѮV��+��B���Q�7���Ȗ��s#�.�E��[
�xFýǲ��#��;���x_���O,�?���j�!�$ts~O͌����9Lu��4�`�N���[=I�P)P��� ��?����l����I:�b�R��kp�`�j�:�,"x�;����vZ��Fw�R4*�<T�1�8�����������i��6��<0�����yĵ}�N������H +_�J&�e?1#�*:ڶΧn�'m�__]
��q����gL���DBbBUU�6IO��3RN5b__m=��k;��.�ײη%0a����gts���=���]��]?����6��o�u���w������-i���Q8]� ���7��>���j��:K�8����*{� ��:�yL����A�$�V6Z���Sv��Ҹ�����|VY���.�}��?�D��bט>}�tv=w�{���#US&W�(����*w�e�Bk�[�������le.ͥ��;�#�u�OR�k�-���TO���f7��V�9��a����M�6�\cbn>>uuu)f"߄�c~���FU�C1�*�ͨ�K�F2ƻ��ر���>�+_�'jЬn�������Î��ȯ �����@#�����Q��qg�|Mۣ���~B��F��\Ğ��~��޿��08 ��j�g/�ڐ:	^��i��+���;5q`E��a�����A�\�$σ�O^�\Q�&���H�;I_����Q�R�Ɯ�Yh(Wz��b�A��M��Q�_^m�Mp)n##M�r�N��c�6Y�m
��5c�M�bb�_��y���HȤ��R� �A�ň-_9�2�G��A^�Mq�����h��n����m�ja/��d��w�a������3]]�T�@1�3�z��V�R�4aĂ��d�"��%�@Ak{X���f6ҫ�����s�R-��±�b��G�KT]M�aW���E�8�Ryͧnb E�;	E6�3�K�Ce�*]�.��X�5����>��
�oj�P�ߝ�zě��m=垕�� �z�"�Jx�<��:i�أ�[Ke�=�~(�~�3����	h��/M����	ȝ�ޚ���{��=��������ׯ_95�u�����"����XfE��v�1ܤ�c��x8���~�38ϵ��ċ�`m�����wŜN��}=���N�5!N��Z��*A'_�����"���2K
.)�N���N�����q�0��ɋ��́���ف|B>���B�X"�}�뛙�圀��(Q	?R�AQ��ˊ:����m붻E�ы��j;�����O{��l�gǸ����x�.��
�c�%�v����R��Lu�q��7E��*��B}���g���Yf��k�����k?����Q��!RF__.�b>\*i�RҨ�F]0����b�I��p_9�_�ǎ'�NO�R{z6T]�^��V�÷�*�'�t���g��K"^��ICZ^1�y]�����<e��.2_U;tF�!{����z�	�_T�E-��������_7��N��A���*s�C8e���X?00���"�;���(�)�!�muaģ�����{y��3����|ċ#�)0������^(��a'7����"5�-�Xt�c	
	����qLy���ɥ�je$H<t��zƸ�b��N܍@?�REM{SFPETg�N�V�x�����|o'�!������0�|���$<Ih{BޱP��]�Z

YY[K&o�S(Ny�Nz��Xi2�>��"���n�<�;l��VX�[*�6��5��?�Ub���)��4�7#�7�s�$�ɠV����oj�AH޾�.b�4�5c�2�����p�s�śt��B<8��$ˬ3��=�A	�&��L�=cW'�m�����᳜!gE�"���H�5;�k���,Qr�
+^��Ѝ���������+������ҖC�THr��%rv�Cq,[���<��,?��v*#<C;ϼz���'����c�`�����'��/@Sμ������hv���s������/�z���\S6)��]M�����wY7��L���*Ϫ��NU[;�˗����Rb3����amC�W��ƭ����7Qv]^��胩N11&] ̍%<�zb|�c'��K2?E9�D���U�C91����.}����N�����l�m|�O�H[6�!�5�~iXf�d��0�����ܽ�uw�;O��ˮe���X��zfK@ qa`��t�t��9qwd�O�Y�O��H�5���(@� �
f�����>���?�jb��"��0�)J��.M�����l}�JI������*y��b�Q��Z����Э���.�����K=fL�ţ����9L�k��Rm87zMH���3r��º&u�Q��$���@��J��-���
���v��N����;k�����x��,��4af�ٗH�>P�&r|)�癦�ZCx��,�1��{��C�v)�`������k�HrnL�To���;Q��>I���ʭE��p_2K=��"�Z�1�Z�ݛνhf�[j�ЬO�sQ���2��_)o�$��D�����1�`���6$�z,�U�a8?�ep5�F����SW�F\�|���VP~~p�"Jm�C��%>�m2��!�sP9{Z*F�U���Y��P�κN��?������5ͯ�&_�Q�?�͖@�\Rեۏc�ۘ~R�$<���v����e���D �JO�J�^W&�q��<F"���A�x*��]��^�����	%�)ͱ���4c]_�p��|���{��u��,WK��`-����x,x����j�Ǽ�\z�C�K�A����JO�����*C����w|�"�ٛ�K�)/=&�۷�Kl݉�u��F�L��距�PT�\�ج��a�Z��Ű��2�C��Ҙ
G]������~d��!�cA�9�M�d������5�T�և:v�+ȭD7�H���Qo�lW��[�΍�L'��.��/�������t��7'������?��t�F���M�ڇ4�+��[V��=�����@��#��6�ӛ�W׭'����U�l�=���� ��0	Ԉ�U�:z��*@۬NM�����U�Ue��J��b�xs��b%wI=,+���
I��c��&v��A3P�0�0�6�83C`�qha�c�Z���Ӧ
���<���B��t��d����njḀ~��Ο��!�*����1�Z#�	꣮s�)��Uܹ,}��~M&���;#nh7J����k M��E~�hɼ>���z�|���ߗdb2���KQ�l�� cj�|_~RS�^�&� ��$2M6h���i�o��H�J�_Z�9�����1B_@�X��i )�@BRP�}�Um��&�9��S�3�1��w�P�]Q�Y^��{�l}5.?�:�1<Ree�����#wJ�X5��T�L� ���Q���a�^'��Ml����`��;{�=L��᢯=XZ1JԤo��c�{]�2y2[V2X���O/ڛ�#�Z.EJ>�R��GWN~�x�̆��Y.sZ]��E������H�h�1#Tw�ۿ������y�e�ګD4�?~�Ww�k���Y%_��	6)���+������}����=9��$��4Q�EH�S�p��ȸ������ܚ�f4�/��ϐ>��q45=~v�и_5da�1�\dQƨ�(_X\��9	��gZ�W�̶xr5�dո��)�B�dl��gUW�H�8��-�b�ijj��V���Lc��������666Gܚ��|�FI�e�<g���F�ll	�Djkj��G�N�		���`�q\?-YɅ=��yD	���>`��&��� �<��S��ō���[�"�����l�c�g�T�՛onn� £Iy
�{;��,�ѫ|.�
5j�!Gx7{n���R39���&r�o��x��i��՜x�Rh3,��,�z�9oگ���6P��wС2-���(2�r�;*B� ��b�V~�{s��1�T����̴B-�aX��ҷ�����[@6�1���r�,oB̍�'+�<�:�H��Kg477�OUjA}�h;� ��c�\
���U�t5��xZ�W�W��(T�}ʃ��!�|[#J�	J0������+O_$��U���W���3��r+���r�RLh=�.��5�E�.����ã��a�`J�oR����#I<-�����ں�x���5�("_�֪d���]���r�Yt�T��ȃH��<���o���㲦s���l���J���̚FV:����:�.��/��j�>�(T^���}��k���r�+��P<��$��f7\���h�����l� Obh˓��C��y�^E��X�W��zd��U�����r�f����֑l���l��`eW0���ASJ�7��9�㕋��|�+�/m�_?7�#��#�yG�B���m��4�-�? !��#�͸�����2� �>���/����]�JqZ����0]��l���l+u�nn�Q��55U�J\����ys׼?=c��⹬�H�Ǽ���C�����i=]i�*���y�="�4�����Nߘ����Doİ��w��j_b]֎`��$�b�
��t�C��m�=᜵�lrL��M`�r�Na%�D{�yRY4 �A���_b���xR�U���Tҿ:�>��5���>;�o��{{&�v����b�`�d��w%y��ajjj�}����}4R%�jԡ�tڥ�L�R���1��I��y4b�>}����pًz��b邝h�'��-@9�=O���Vj�J��Z���Rj�L<�����m.�s�A�X�0?�	�y��#�V�����v��f����!�D�
��}Z��"��Q�VrQ�C8�n��?��(���j�	(*F��s�ұ�ԫ<���2=+/;�!��9����>��
p�p���7+�G1��iW�l�l����U�l����#�j��a=�WoS�Dx�t�#�
g;��[��7��Z>�ڿ��m��b���mM�)��?w�,:+�ۢ�+�����������|�t��~����rD�ʤ,�k1u��\W6+����+B5��TP#b'�9�j�=�;h����h�
�:z���[q���^�w����N�kq)R��C)����������s.��M&���L6sYy�z�k�`��:ƨj"�艄?��[+�⁕���b�& xޓ�������+ʅ�d��x�
()Ȉ���Ђ�6<h�5��]�"��Eо��<����U����`�`*_�!�~_ɩE?�	B���xv(�F���O������?u���4�����7����Y�_��(z�)���S��DJi�,}_��_��cW�
�R9p
6C�_�;�ʂY��q5.I�/;�j���W��hR�Q�4�g�i~=i���*�\��D���%��cv'�ʤֻ���e�C�7_���^e������TR��BX����7~vvF��"PZRXn���V�|�}>-B*bo^;�;�_���2݅ʦnQ�xt:]׹�L[���V��[KU�c��86���i����m�@;��X�i�[�b������%��QwEEE�]�i~���'f�	Ӵ����	l�?ߴ300d^��UbU�)B<�R+|�_l|�c@��nߒ��m;(0�y��e��������ڛt��3���g�uv3��w���:�������ڌ/a|=�i�Q}{���z�Ux��G��־!�g��h���/ hL�_9��>�7)_}4+�F�����_:�Ur=�*�{Z��d65=="WWD�=�&�����lA��oZ�<̝�ԉ+F�F����V)��n��W�U�r+�)
������k���2Ӎ%�!�̥v�M�g��/�[�XP�hz~�_����x[W�>Lg�vW͚���t�\��"�X�)��5GVʝ(��2��RO����:�(��l��1l��{0����A����9��-�z��ݒ�b�Իa_O�s
��P�0:�z��#@�\yc(��
��=F<d8��Z�����ڨ�6%	u����L/���su`����Hs֨�i��R&mt/�oֿ^����]�`h�QUO#�!����X��]� ~9��]��TL::b�����S�
�9����JL�(P:�}������aa��'7��4��j�'PWo�_Gy�k"����� �qyg�������`z&��)��娕
�b3��{�t���9�Ї��Z��c��j=h�		񳚌8� �r^����!��CZ&����*���zh!��@��<3r�18�qa�\��6�U��������~���r���	:���ib���1?$�/@j@���+���T�h`沄,�������� {���{z$C���U02����\��
?�)�/~��Ⱦ[��m��hO��T�I|��������H:���	o>F�|�8��mO�J���l
������*;��k�6=�E�I?m
��5F�/�ִ%Y��f*����q�Kv���mY��9�dB��~9�� ��xQص(���2Mq�ԧV���dma�҂���3Q�3�"x�-��y>�p�j��7d+>��z�����&�D��� �zC!��w����E)�_�;�����6Cq�?����
:�$O��]q�0��������G/�����*�Ñk�LT�9.������X����ko�v�ZW�"��ii޺t&vh7�~y�[�3`^%n�o���������2�:N�CeY�r�;���p�/wg�#�B��_��U�v#i�����m]��כ�t%�eaA��IPĒ�AAc�DD&� 	�� xz6�}}`:%P��RmV\��+	v�/,�S�/?�Tome�P������W��ڇ� ڮ~l����-��y*��|�(��>� �Cʏ ��CRc���y�Ӵ�2����U6g�5w�N��&P6v|�q��7�-����:t�b�4%���f/K�d�x��D�]c��+�0K�$aA��Mk{���?�-�z����e!|ԛ��'"VKC~�K_cK�'%���G?$�QT�ɭ��r�М�92^�j[^yU�տ2
[U\�O��)Zڔ��M��س��!�1J��$ʕ�㭖����H�»F\�<A�+=� ��e�H�#k_���U f�*�!`gBǫ�D?C'A���̇���o>m�Y�R�<Y��:���_��Gp�@!8�Bo�O5�U�����d��c��@�B<��uɐKt�]�O��։}�0�j�E�\��2��-~~w� �B9��uҌ_oxf׶b�IЊ�w��f�$���X��pI���V`z�芝��_�������C��[������a���	�ށ���"�%��:ӻߒ��,*↸��;'K�P�zT�%v���z�������|&�&��u�w�|��S�X;9H.
�����(k�&RYY+P��^9�D��݆��-(���:#����T;�H({D��/�	x��ǜ��l������	gZ�]�\L���h���Uzu��'`)�Ć������W�T�ԆR[�TEP�N����������~k�AX%�B�3�>F0�x�� C�'	�����	LX�-�?��K��� �O\���� E�����`��i߃�0��@�%?_�c�0"V<-A�V6����!&]�Ht�`���O�mc�5ߣ2�����_C��S��MZt]d��dʿ2��l� ��З�ޯ9�|%����#���BdA��P�Uq}!IZ�����U�%)�h���
��}O���(�0��y6��ڜb�y�Ì�!���IC�,
����>K�ql�ͦ���t.��E:U�i���,�l@����!X���$έD�%L��H���hd�Ȳ5�a7�\$�x���d+��O��Hhʦ%�<o	��6E� ��X~����Un�h��ѡ���
J��>ŭE@��gl�t$6����)b1i{@�p�^�c�#�M��J%Z,���x������q��Kh��-�'�$F�Z�g�YOt���|�i󏊇�{��	��6ҍl��O�m��!㳳c�����hV8�bIHN���3l��.�N�X-�G6�p�ТU�v^��ػMfI� ���L��	��/�m#G����uc��x��9�L��A��h���=7��7��\�}�$t�08�PϦbV+�v���\��˯��p̿��!j���Qi���Rؗ�P�E���q����(Y�^��D�ä���U-�L�J���{��D�Ǳ��oxQ���p2�Pc�iEh���	�{w�M���x��s��w�4���Ə���Y�;�#��ӱ2��ן�� ��H2�K!�73�bC}{XU�{�
�P�����gͩ�1��������GF;Y�r+�"Xm͇�;�腂oR_�����t�K��L�I�E,�
�w�x{܏OM�pZ�O��Z��)+fuy55跷�66HF�C�t\��<�.*g�>F��VX�/�[e�K;���4��$��ق=������`�O�1C׭�U�����}��{�|��pB{���ۣ��D�Q>Scf?/GW�z��(gEc�%���G�2�ϸ2�"~��hGȨ��u�_$}d&V�L�kC�����w�ץIL�����4��u�^i�$�]i�bz��"��Q�iy��Z��u9lTq�p|�r��'-���Xɥ��`���)��Z��3�|*��hPi�f�ܽ�n��!��&�z�,	�ǧ�/���i3:1���S>=?��bo�ΟT;���j���)��||3��&�����O�|p��,[�O%UT03��Ӽ$��2]�M �	���|9g#}�Z7kE�U��OՉc��7�q}���/�|�+w����#��s��q�\�Oݼ���i�p��cX��3C ��:��M�������S��B�?��yW�V�[�Sr�����}0�:��>p����.�qo�@�6��n6�Ɠ(�_�|�Fi�GY��Lc2�N�������٘�k7�$v��wv�mv����_3�<���UUB�R�#`2��?�ifx�����e�Az�����)�u*��m�"�f�rfC#(=�;�yJ+�����`Gj��w=���x�
�S���f�Hu���,���:���a�6C��?�?�skD�Q �޼x��kh3 �Sl.C,\�.�@���Ɔ�΢�D��vp�Vp^<���:"!?��[8+d\	��vM�E��� n��᫠��D�ڂڒ2�(�E���z|Nv�.&�"ъ�wo.����J�&ۭG��o�����g��R�^I�X��G9B��Vi69�����O����3�]@89;\��l�O��@�vERV�?�O�oY�~wBN$d��������8n����E��f�D��U�������3U���i���\�>�)������6����]3���v�رL�`����0m��[��ɘ�0�a��޸P���J�T^��}�y�� j�Z�8�_��Z9�]��]�j�)�:[M6�a����vF���![���B�_X g����ť�Ww��e〶�ǲVN�G�^��E_<V������_<@;+=�(��λ+tT�n���y�d���*,o���6Df_D���޾� ��������-��=�>����{�iz�����<���0�b��e�v�t��\)�ru�N�Dx�T&	��k'g�B���xb>�Y 4��ﲗm�����P>�?\	��^����@��<��ZԘl�b�Kk<0տ��Ɨ��g��^E�2���L�@�`�~��g�;��/5[D͹`��SA�r4k�ڕq�1�M7�m]'��hEb�"I�Dn�n�a�'��+'�A3�E?��6Ju?���]�l��k��t���Q[ʘN�.ByӮ(�����c�ʸЅ�W�n̸�/� =BL}\���j\j�Y�Ђ�r{�������K��X�z�����
�U��'(&{$_@F���\��<��U��F�W�S���E��~!M�� 	�~�Fa��m�B���"��%��I�������L���7ůxُ~�`a5���J^��RE�]I��|��e91'��:s0����5�NmՉ��^c,`�����_|�U��?����IBml�jv|e|{Z-�<C��H����Cx��~�^)��'آQ���֋�"NUG@��?7�����
��r��=\���q�s�6�s������������W�&=C<�{����_{�m�vTGf�T�g?�ѳ����D_8o�Vq��n����b����=��N�4�^q�E������8����l�,�|VE1�XT�2�Ս���|�B��b4���"x�c�M�U�K��dH�	�9��1rå����.q����������jKt'��W��� ����f���R����2�)V�n;Ѡ���8q�I�j�_^��n1���m��Z�)��9{	�����������_d�+������Ӗ(ۚ�r�^�f)����	�V#kMr%�?��������אE�lV짲(pU���x�>ߛ�ee����
��\]_ǧ�G�ܸ���?�Xse�������+jjFH��������Z��SH�������,���L�Y�SL.,D��,7�>ߟK���Dٵ]�U�?�=�����l�����Ԅ{<W���"����5�J�#�EB�&h��� 
�=�9���CI�������S�m������)v&dWM��n�i�9a�[�����#���W����XW>�����;��z���C{���U��P���N0,�@��6�Æ���:	L�͉) �DRGv�NjG��v���zt���C�v�}�^aK4�׾<m\7~���U�������'��Y �S�a�ǔ�V�A����58�\
C�R=�yY�V}�/d���Y��c���̅��-U�!n ,~*/
c���T�S\6⭏�<@N�����MxA�Ŏ�&�FߴN��5��P!�_+����絥X�I9�1Ǉ�=�3oa���up�3�ܟ��$,h��c]�a*i�C]��J|C0b�GJ�G�I�0ɂn��P��#�
�i��~�4(]2����j@�;;���ޜ�d7�zw{��#�\�v�X(;;���lZZ?��l�s���e8Y@M3����I���^�=�]o~y�Yq�����(��**�^8u�����᧡�Uz,ܩ}��r:Y�������� @砣b�jDd��z�o|||`w0�;����h��� ��)o�_���ق�����x��aXYY�7��';��s�|5��\�"[e&�9����n3�j����c�@;�AJ<�s�z==v<O���m� ���#�;%]f� �g��]o��J}񧻶�����۪����c�����\�^tP6v^G��ʚz�.�د��ˋ^�g�}X®��%EE�	�+NPJ���g����B��|	����þ��{a���T��.\�4O�.�	��ݔ�1�S����;�	��B�o�ݣ#+�zj��dY�����^,�G����m��2��D*�鎅����)N��&,�b=rϿí�����
Z�������K���qq.,���zj����D#���퉍MLڗԫ����K��l��[�v=V�Ym�֮x�ZZaʆ���/�}�mog7 �Uho��{ӆٙ���G�!7IYY�l�=���� �@�4|����%r�.�i��Br���0�~��)2��q:��.����:���
�ۗ#�GG\�F�F��hҘ��p��3:��4&�|������^�e����Y�,�Fa�v��|j�<�j��zo�z��)�\��? �ZPf}���K��U�ZSx.���l��L��>�˧(��d�7SK�B�Ow	&'�I^3� v��_�>�q_�
�t�M}	Td5PT�/f��~����i/þ���*@�h$$�!!PU�e����{/=Ϫ:����a(��Qx��`W�]c1�oG�	��8�ߺj�-��s6�~�c|M�`lAW5�l��c����_��x��y�Z�}������0�� }ɳ�$��:ZN�iyǣ���c4�߸LǏ�A�^�Z��P���_��ߔ|���[��L���~ՌȏH�u3��P���<�Ǒ\YE�}I>�'��H�D�mj�����B��K__��~t~ĸ���8�L�L��F0�t �=��iOjh�xd�mt�O��Tƻ�q�-����{ �j�0<8�;���sc�קb���b"��X'Z:��V��ظᵵ�-�۽]Z�)��y�#�k�j�<����	<�rvC�o����Ε�Q����I�[��W1Ry*�(c��Pdk>:Jg�&��A��y��e���p|�ug������F���h�g�^�qgMMw��Ƹ0uR;۝�k��kޜ�) @��n�������������Y���ǀ_�//g ��X;�e�F���ʒ�.L��]���"�R�%;��'e��S��v��(`8Ő$6����'�/s�G�e�e�ᨿ����mc��������6z�'s��
����/�IU����	?܇q�/�B��z��������7�����%6V]q;<�1���j�n���� �);�����s	�)�ݏJ�D`J] �TZ[p��������d���������`HKːy-m@PV����G	8�A��p/I��ɹ�^env�h��֯����� ����rی��,.���-)0��L�EDG�M�;;��q|y��6%6ǅ�^q���x���3����A���s�eAR��>�� ���t���0ċ�H��B��8S���g;	�bk��	Q���y�O�à��v��tw�Y~����c����1AG���k�- 63�J>����R��s.ۿ�P�J�[2P������&�X�j��V�a����n;ٵ�O����egHZ�2~〰6�m�P߮�wI( L5�0�%0e� R������`�F��|RrS �_&�q��� ���Nk�1U54(X/��
��͍g�eL���s����@Q��8)	�A�l{����3?��0"~��h掮x
)�)�������{��O��N{�����?]eZ(�͂���  (a�)�Z4{���N�or�Y��1EK_��|�K�!�dQ�P��H�UҤfw�H;F'UF�y��d���`W�Ҍ.��6V���a�m%����V5.3҅YW�Ճ}��n+��}�<љ���s^}w�[e}����up���L=�<�X��3'�G�Uh���8|g�����IN�Y�B�Q;�"#�2F\�U�=� ��掇�cWuu;��VC����[�iiE�W�a��R�|�7�6ĘL"��n������9�	lY�����H
��o�X���lD��b���U�b��S�/h,~a�&���~n3���9������z�~w��#E˲^5(n��K���}2��˥L����v{�/:�֤�d�(WR��*�y��@bW� �%X�Hd�=��J�g����v˽~���{�Q� 'E�y�`�\~kS���)8_/����n��ۺC�+�='<�,Q��
�Y��1�T�|���D�1� �d��s{���~��ײ/cJ��Gv#+'W��S�_?���V{ڲAF<���kT��m�����A�7==��?�{#�]K��ND�U�D�j ��,�#p����{S�+���B���+Y6�&��F���}3����ݳrf���m'\�$�Bz7z7s���R�7ښ��� �/�T�t
�FV��s$W��y�h�ޟ�BR�l�}ʻו���9#B	2؏S��^��r�g�2k;�|�ޯ�G����WW���/}�K��rx���Kzn��e�k���Ͽ�**/2����wc%���d��}��r+$i\��c�^s>���C�o����Ü�����m���sT��٘L��6��� ��^? ��5���s�u\�+�e�6$\=ޮ�e�uܾ��N!J5��|��(��Z	�����?���C�=^o�=v�X�N4�&X�n,���Q�Ĵ��p�5&�\4�,b�\��e�[��د	�z��GhqJ+�`Nף���C���
EID�@׫��r���4B�8�/�~͛�j�'���֋�����#v��`����M���k"U0N4ܽ�M0\!��)+p������&����E�v������oo��7�{���j��rڂg�7e�
vp��5�ƫ����4rzf�y�'���'f6݌��/N�s
���Aэ�ε�R�c��*�aG�%s�H�����mu�7���.'��Q��jpqn0������7�h��~�v��L�ς���r�z��~# ��N�,`u��@Y��>a�`�x��5{�F�
�Y$�=>�ofUX�	ɗ��0_Y�d��L�UPV'���R����	��
�`	����>�G�F-�iC}��w��u�GrҊ&:I�]�g�Ѻ&2\�N�/�Sq��Q�^��'���l� �����*0X[[�L�;o�hr��,*X�ΰ��{O����:��#�B� � ���J|��e5C�9�PN�T����A�{��u�w_��sz�ԑ<�2�vS4(� ���0#��1
g=���z�-�[H�7*�����6���R�":��'ݥ0�^��ho���W��c�z����*E�
s	���3�mb��:�0�f�|�Q<�L{d�D��T�����t1�/��3���=Q�k"�E2F���H3��חS>w�at�d�0���3�Q#��E��T��m�/�����l�סWM���|*i|"Ѭn�M�pa������z��٨�hB�N�_�L�=^i�6�U�n�����:#�c�O�lB�J��g����0��;�%�Z�h��#ҹn$< �'i����y��D�G��m���@��Fđ��9����Ź
ڡ=@`�Ҕ�d\��h�:d���('�{W� zض$��r�O��8e��EVR�,�Be�ՠ{��Q��c8^y's3�F.�M5V\�C,_�`֠�m�օ�E� K%!��w��?!^����³�����G�u� o
�v�����c��76=�җ��Y���_���Dz^��Q �@�ÿ��{[�<9�z���+�>��ax�8���|�Ȋ�
.�z$�:�!��J�p�і��]�7��9��@����'�����E6P� ��w��%c4� pnA(�o%V��g�д��^�ݫ^C�̬h�������q�*գ�v�7�y۵���١��П�۽u�oY��w'GՂ=j�WL(&3&��/�?�~��@#�b&g�gM���l6	�D�lv
��%"�tvr����lq_���A�U�)�^|B�O�h�^7Ei�" �Yޯ_����$P���l��2�������{ö�z����A)���漁?���I /�f�\�:��9�ґ�W�5���/���n	���"Y�ٝM�E�fҤC��)A�2�5'ҭ&��g�3� �"���#B��.�������,ų�c���������j�
�<������w��'� M����C%o?��<�l��y	�ˊK��k
���ґ�݅sy�v���]��0Nt���UC�����Vqc��;��.�����=�Un_�r�x����pO����ëJ��[��Q��
ho��S��5��Z/��W�.�4Cϔ�٪��9����)+oM�M&� ����|P��]�%��h��|֒Ŋ�Cz�G����ܔ�M�R"���ڙ�C]x^� �1��ڑ�J���U�Fa��ce1KC1�9�+�Xň�{��X�.LR�I"E�y��x��V��Ϟ�D���߉E���_���2p7r��cy*P���J��#^���4��w���/L���9h�r����:KG�JMA�
���r驩���Gخ�׏vӀ#�: :�|M>x��v�~��/hn�󝲪o:�;���W/��xA?T7=��9�i��-{_#��
O�<W��b{�d��#�LdZ�q�sU�YQ����N�'~A��]<�����A^������l���Q��s�B�`!��7�l�5��͍�]����~\;qO1U\����kݦ�b��x� O�&�k��2��A��)���IC�D�Z?m��駃�
���3*M��<t
��ۢ
���A�M�GDͥ�*Z[-1:5�!�����?�+j.����M���ZD��¡f���������EDZoz2����|�oww��h���c�l�����r����;�wH#��nD'�S`��Y�Y����Y$��?�c���X�E����]:m����ȣ�?����S+5;���#têx���a��~zczP�>-�{��o�REk"�k绮��q���H���J|N�(D�*:h` �>�]xC���ͫ����u���;Y���E���'�z�l�!YH��a>�.��wUV�0e�R�^�yw6?7���e��|�����1��x>�á����oU�{�a(c��fz�M]�Yd�_�ߐFl7��~mlNiv����$/,�R�gB{"��E��o|'1��W��&��
\Z�+P���F(��Z-Tە�um7��|?��)���?Ӷ�U�-�j��{�U�Xm��]�5�z8;+.R���[���*�؏*EK�Ƞ���E��E�ɻ��hͤE`�z���[�oE�W^���%�C���]�G
�E	 LHP��;u�s�7[�8pb(�]:��Azb��<�_0-�ߐ�9����r�y3��=�<p%>z�#t&>v��[�\�/3��8����YFQB	�Rm\l[��*�����qC����ìz�zW�[`f(�� �$2���	�9.L�B�b�֟ӳ$gB��+ҹ���ލ��a��@
O�}�1x�w�B͘v�M�8���,���!��ޞ�o������`�M��>xB^���ӣ�*���P��A�z;�n/�(�o�$B'��y�Sr���ʠ����=B(�d:++�b�j�?��-������ ��5)[G�G�r��� k�:HtU��Eԫ���`���LRNH�6�Ҍo��]�^Y�#�EV�Ox���ڣD���b�yB�H�L��ە�I8݈��[��`�Y������>.���X��V�@PI2�t��!^����K��o�����\mu�K:�#�9	mN�e= ���~:XD���fݘp��b?��n����������ߖ�4��Z8�����圎}�v�Ωb���ġKDt��ϟ�f�8Mkϒ[�%c�z��3
㠣���L���y�N�����������i�5=t<z�,\��<�������o[R���a_*4�b����}z�-�ڧK���[+Ե���2����u�!X}�1l��i����;���\gv��!q���d�d�m�;Mɉ�g�,��^BB����b���u��p�/^������!))�ˬ�۬.�E��w���A�m��E��'u�[�$�}����R�^��;N�lll��;$!�O�(���4}�
.+AA����ږA�ggǴ���5�n3���}%��Ħ�B�qpч鮮����_�=�xbz�Q�" ���Fq>U^�ċ����VXc��}����k�L���$�s���r�`\���C|f,�O�J�#=������l� ��*����	�g��³$�޹ph����yEE�X5C��7�����>�tG%��l�Ƈ �NxQhH�P+�h���Hh����1{[�Tbǝ`�AТY�.�͒-d��gD��� ��:#��%�k�F�$)�����d<�֍�vB��@)�Ԧ�:S��e�OG��w׈�AYp��~��x�{���~��NDddw�L'ME�+��!R1;É՚,�HCcc����gJ����܂__�K���8ݫw�cR����KJJ����»E|��}wrғB���_.�����߀Sn)���-��I�y��1
�Re2X۷�	��J�:�B	�9�U>#I���e��mL�C��r�nXܾ�s$�=֑��
��vB�W�+����j;�P�q�C�[�'q�=�����F���w!_Z���� �|N$0�H��Ƅ�}>g�a�>��Z�@�v}�8� �n��i������b��R� �Ӄ�o�:�H�B��)����}�7�q�Ejc�����#jjJ�o�0�U�}
O�z48$=����䳝7��Q��Ӏ�����\Hr�-���C+K/�3/zؼH/�Xv{S`\ɡ^�����$d�պ��ռ��2~6I?��O$�z<�R�I����qS��m����V*7�nփ��9�����f�1�z�f�Ã���9$���B��i��O�}�\���睱��s�����
OKK�tm]��/�kLcr���Zk\��O��vvv�ϙТ]w��5��Q(u�Q� �sI���X�%#lAs�OǶY��P����|`�BGI�.+1��?����#�
�V�pd���/ڕ=�'&�w�A�wPtl���A3|�ec��]��4�t�'1Svx�{�p�ڣ���x����I��a;Z�NVQ�F6�jl��WX�j�=�H|� ��}��W�N��x?�o���9�#�>[|�	A����ff��Рf
�I��NY"3O2^~Q`cc{l�蟩�9;;fii���ZW�uK��@�`��wk�8gǺ{�ў,0)�)�ȩ����U`*JK���qAʐ2�4[ZQ��;r��}N�������/��e�ʥ!�-$���+ikG���3u���-��Cb��
�����D��ˎUum�ݞ����#+5m�F�Xd�6),�Ў��� j�2t�|��⡖�6�m���4{#�		%��H�2�V�0#nw��,_��D��?iٜ���Ȗ0Ƀ���rΚH�LL����re�c���{�!Ƹ�w8�0� r�.aM�#`��C����h�g������Ta�-���&8i�r��-���s��2��Ѕ6K=`u7d�(|�0$�+�UJ����љ���8�J��C]�[&�k�/����晼"V&��}�3��UE��!�y㼭T?������&׭�y{Y�hM����d�|Qa��f������}J\ř`�܍��2r���9����(��>��KJ�5y���&	�k�cL���QX ו�IR�*(�n���$w�Qt7���z��$���D��0�a�*���_��W�o�C0�O��T,v�C�+h��{�:4�E��~K��Y��	?�Ʀy,��e�}�Ӹ�/a'�MƘ�MN���r�ݦ�i�Ԝx�L��w����tFrb׹�i�
b�9������
����iP��x�|7�$���}	��� s3���L�(Ě�ڑy��z��ߋD9��r�p���k�2�W><]3��0=����Ͻ Z���fb��pZ4q� R�8%(\C<�����B'y�t9�(�� �<���0�� Z"�?[D`cg`Y�j��vt�ɖS��6� ��d`=Q�z������BK|��M�Eo���0�"(#���c=���
ۤT�3a���!ˊ��"[Z%���ގd~�557�S����Ԫʋ����݇�N*g�O�8�-�Or�W:N�û�#Ɋ�X�L�f`��VI�3:�,��B�������t�3'�#�;�l��lP��E�;�;�5�þ��D�pv+pz��d�=���K`��>�����#�va<�ZD��6ıi��E����'q3�G���M_I;M5g
��v�Z0�S����g���p�s��zl>3WIYd��.��A��+��6L�sA�����/ɺU��i�>��UԺ��E#�^���䉏j~4~��ڡ�)�U��L�DH#"Ip3^�c%�����̝{6t��d��$��h�����5���ܑV�z�[kDMH��t]�mb�H�����)�Sߟ��Z;�ʑ��:�����M7�"E�_��x��ԋo�U:�W��K
��83����$��O�����yRB!�:�=��y��̂huŕB�-Á+s�P�2W��
IɎS�@_��RY��QCOگ�'��t6g��ƂOD�U�I�М�u#����{�ڈ�<�YNÅ4�Z����Z���"�S�	q�_P+�U��Y��]�}�����m{>�HL�G�K��ۀb%���R�#/X�������ȉ���*,����Z=!�`ie�?�� �b-i�B+P��M`:`C�p��X�(i��P�8�
�8���IC� ��Y=D�wL�{�":�I�����K��V�K��  �6�󜹥p}hUO�8��]~]ŭ��܌�_���z�e*��}��CrD3�r槲MIT���ǭ�������L�2U�򇯾���S���2F�Mu��-����6��f�l-I�Myl킔� �±et��\bsP+i��%���=��u q�7������x�1�}�o�Ʊ����*3���훢5;�-�Z��wq�1'n�Y/��K��7�0�s:	I�j ǆx�.57�Z��"�Md8��S�b��x��"��yK$&�j��'ݍބ���w �����V�_bY$G�d���~wR�����{��3�6�sU?�7�V݁@���rEn�=>+��X݈��_}�[V��k�/�T99ŊU{
'e���G���s��a{��<ιdg#�V3�䏠H�:��Vч�V�y��P���5̨�Y�ߺD�t؟�,�5%S�D6�����!p����O�ש��M�z�ϒ��IF:~����K�\��Hh�u� >Q�@����}��S�@LG�g��9u?&�r�i7{�n�9S�@YE[1��#��R�d�kxP{��n��M�Bϙ����Q�����F
{������J�__��,��%��\�5[C���4�M�M�]q����&Z�?g2����$=�ǰ�D��T��F����C(S�̯���y}��[SqӼ��x���^�����[]'H��7�G2�l��ƺ%�pH��w�o<*H[&�y�33!	���k��[ϻd��i����j�/�������h�|�&q���^�\�qc>�����*�+�A�s�ח��.��Am"�B,�z�aJ��cʇCʛ��L�@ހR�S�HVw��.�����p�Q=��/�����k�zS��4��h��	,x�t���I/�AŁ����7������ΕO�&mRa��a���F��ε�~�0G���7mH}�����joƚ�-`�uΊU�Tx
�~���~���ȱ�_.��J�+z���2�̭��{����D�5���}~l���+��(B��i6��|z��O�s��k��c�!����3H�/a��X��	�oR��������nu}�{�.c��ۋ���T��an�CڂՆ�i�[Z����l:�����&�ׅ7�:�� ��y<�W��T��gV�`��/�����L�Y,�&�V[9��2s���(��;h�_��D�0H`�αP.��(Lu��rN�˵��;������8:C��'b��	/-�@��1�M�pg��J�yN,���-5C"��񘲥N�dεw�n{?�������;�)��ѐ�/�
�7B�%�nȓs�C!���&�R�;I��6�*]�z$W��Q����
R�4|�(L�2r����̐�JUu��#�8�]��D7<�p��6p��p����8N����"F��3���������|���vR���vg+H���݆Ӈ!��̓��Zk6���Jt�f�^ ��9�>UN\�o��F��k��
���+���̵��$W�؉����^I$���q{ߡ�_��r�(��`�G��yBQ����m�?�0�+(7��0 �ڏ��:���sA�������I�.�LMA�;�,B"k�j%�n��8xs���̏4�w�Ӂp=�ߡ4�P��X-&f|JJ�&��1��Am8���-X�"AK�R$xpw��Z�xq��R����Cq���)�/���ͼ3�C&�{kϳ�waﴲ��yn�
x�8/�ES�<!55���!�O��6L\�CQ� :v������(��o%�zǌ���׾�������^��؃���r[Z`
Lh!_q�&�cb[�*�Q�}��v�+)G�7��hbi7���v?O�R�raټM���5�#�F�O���Ҫˀ�ϼ����~�y{6��?k�E���fu�.��/O�;Cy�ؿ&����_�W��������t�>j	�<jB
PF7I�سɔȘ����J��D�-��&�9����8�ڢ��z#� L x����F�R�t�똯�sR�s.��l>{hG��G�P�{�_��>����(�	���|���M~���n������� ����&���h8�c����{��G��\M>#9��c����0�d���Thy�7Q2---�7�c�#N��:�p���]4پ��laVޝ��hɰ�r�NȎ~��5���;���sv�fN����5���W('��}�>���>��� "S��k��_����=�YҖ��}%�?c������FW�ۛ1V�թ���Ox�t�٣G�J��Sj%�o���s����ǪE�"+ѳ=:մ4^�&�<������������l���|=T�����p���ɪ����%����Ȓ�Z2[��` ^Kw�<]��Q�?9�˛�ȓx�y�6B�~A���h�\�k����a-��-u���Lw�i��;Nȅ;�>1�ݮLI�O��"Z��	��#l!�������>�@)y��?��4��+>�3K!�LL]!ӎ��t�t�?m�;!	x�_E$�r�v�#��z*�b�ڐ���'hc�ρ�+��|���8�;w�4�M��288;�){�����pE��z�hR�,�z�Lr�A�A��4+�T�u��������]Z�#�������A�h%S8۵��q�(\��Y􇒁曉I��F�3oּ��O�r9Kb��J@�f������D�/�~��J��h"A�/�À �u(���qqY��|~>���JAVV�ʊ��7�����3�l�c���7F�>
M]��@�猀\b���lEZ��V||��Ke�V�jB�d�i���9C2�Ć���_ҋ�0,�x��@��*��&�{ L$:����{��$�/^��s��\Z���X��-i���㯆J}�Q�2�m%mkOTQ�0�����)�wg��������̙�����֩e.l���NXMEi�sf,��j��aXV���K����l[G6jAO���޴��g�ՏиӬ���-[$�:��3!�<��6�($�L���-��w�c_�;,2��c/K�,�G[�~�0��(_�s�3���fv~>�K��6�+a��k�v�}Rb$����̼�+�I	)`_RA><�u�	x��E��w�#������֯9r�;rO���vu	��mnm������	���\�tX���b�����a�3fR{E��a�`�I=8�u��h-�z>�;�6gPs�"�f0��BD��v��޸��$����k��mGLՊ����A�������c�y����U�D�U'{S���~���e?^�^�"��@{��A�P��#��7�+��ܩ��\r��S�Ϛ0��������K�HȏV�V-Vh` �;L�sZZ�~>�y:��Y/1��������"��6��f8���_��]K�yˑ��[��`ەs��OJ���蕈�	�pT�*~������EAӾ�y�4ԙ?���L��W����E���
fL��r[��8�=M]#H�4k�
g��yKn��`����Pp�]ZW����S�c��G���400�?0pF_/��^	it�K-���d��~gmrMD;a��?@���k�MM%jzXTQQ	xU/�ω;����e���1�%*]��ޚ�[�4O~�_���=�Evds������&����:�i���?�F�%YS;�ڑv��!N	�e��[ͳVu]G�z]+ܮ�BU���s+��UI��	�x�C�cN����0�L^�Q��!�ޝ�J�G��bzz�5Z{�+ߓ�C(D���@�̷y����v<2��^<x%�fN�2�q����Ml�[v��s��C�"X�0�,��v��@�2�JїTؽ��b�3vL ��B�I�di7��q��P�V.���j��5��<����6q����dN���(O�����[�X��o���49`��^���K	rx��D��;1
z�]��s�P�s���i�Λd�{>r!�̴�dé^�Ǡ�W��	=m��+�M�ys��7[��L+��*���V	�(�ￛ�f��|�0{�l�O��������e��GfD���
n���ߕ�@���a'u���NNAY�ލ��+��XO	2�o���3��֥�$����|�"m "�_��U���qU]*7���	�?��~A�U�Gզ�c�nA��$?��'~7���PI^�b�.��OL����f
p�]����wR�q��w^��=͆8�C���:��<B������DOm���NξaPJW�ي>|�,Q��a�:��㸽u�BՑ��7�����N��4AQCH���/@R^H�.�P����K�"
a}OJ�nn��D���w
���`:(�FTSS�k����к��K�̯����t�s@�`�OېI8�?pZ{��0�.�16O���+H��.	�Rq�P��!�Qf�H:
��EN��{΀���O��ɫe��G��͔�ڟ�	^mY!
��<�ZeW)��;��3�^�g�y��K��+c|y������Tif���a��/��H�����6����I�4F�w��˔�/�o]��o��W�	C~��v��O�h��{�9fQ7�H�=_�O�8�Q���8�L�|�Ƃ,��2����bB�6����#��[o}\)FV
�1�ơ~��V�*oH�v/�D���){%`�ɝ�n˲�49�溔��`(���Eɺ���C��������j�"�6S�B�npN����&�)y��(�z�oM�."�47	#}K}�@� �A0r�p���)l�q�y��T�_XzD8X�o�z��pZ��ջ�+��d���%��P��F(�N�	����[D��sq�������9$7�����9�:F�)f�bdymu�����#�J��z���r{QN�]W�b�8���jE�W�0�zN���ƉW6�/J9���XG���L�t�ε@��� �g�h��Q<���-&��i����|��iQ*4Ƭ��[k�7��i"�f��-i�c췡��y};$��&���.�s*]]�n&&&��	l�;�&�����_j�/�;�5��b8������"��!a�M��9�$��͌2� i� f�Wz��O
&�a,�
���'Ӱ#s�⏰�w�E��^�m0��uB�	���,�c	��d��Z	
}8l̒�����������~��0#�Rf�7��m(+��R�p}��oCq�ݮ�N�kD_/\�f��j}�]]�#���|'���Ym�[���8j��&���]E}�שG��f��F�ܓ�B�kl��9������EJY��^{��@�"���j	�?@K|8WQ�:l s#���$ �Diώ��� X��X�2:)��4�.�2%�9�[��>$��p!�@=����$\}�:�%-��JzN�G�.�=��]���[�ѥ2�����,��>3�`h���d!��B��,��+�y'��RZ�u U��LȂ���S �pf`���\���A�V��E)��J�9�h�U�P��8�5<����l�y��%C��aa}��=�C1!AB�0������8��I��I4�a���Q}]-vw-'A�c���CM4v��Y�f������Ͷ;si����/G�ga��� &�Vσǽ������0�2pa�?}z�K�	�2>C�h�s���B��P?�z�����7Mo S1w�_)�`k�x���T� m<��+%���I�ƕ��\��j7:�	��Y�]^%<��`� I���m�Nm����`�h�jQػ���I}����>He�Uo766N��)���A�[Z�^�̰g�YV8��<.6��n�-H�E	
6������$�i��B��I���r��wy9��]I�_c;�!Y��[y�<��"���?##CJ�����A_��qz�h�Lڴls��.P|`
����۫e�J�� �6~C����9������(hs�Ɖ(s�e�c�H@ 𷗕����Bl���7��h:��F0}��E��^9��ճ�͍tC�TρZ,���D�Î|`��f:�1"**�w"�!~Iҩy������BH%�YZ���F�+���c���KK�Y?j�7`P�jK'��U:�_��|#�1򎎨Z%᪂��X�PvA��R&Ћ'���bF=r�CQm�Q�[b=.���+���v�8��;���A�t����242�m�$x,M���L��q�pWr��W:�q�����H��1�Oj���m%���Z�Ct�&�MP��!���f����q��SDy�4�������$��u� 8m�C#�I`nm-w�N�!����V������&�јV`�>Q��7(�F`L����L��e���z��?;˙�ܦ�	]f�Ԟ�����X�����J~��`�	4b��>Z�A�(������0��VO)�a.6��`[|�"E蓆��GVr�Q8L�����TB���;(N5ؽ�9fH'y����`�R5��?*�{#�! �a��A�{|4�����]�q�L�d��ڰ��YЅ��X,��wl����`�����0�3�� �6K�B�z�}�:K�S�t��?�s�)VX�98/r�k�U�є�T�,y#*����@%���35�Ľ.+�$�8��������E�<B�o�	Φ%�7JKҜ�.�j���g��̭J|��+?�v�+���2�B.���n���y�
�%A����h;7SHM�H}LD܍�v_�1��z��fo�4�$Vh_�N;n ����^y��e���cP3+_i\928�<���EA!/�9_�n�Utz6.�?��1�2$����O�����BJ�Lf�YCDO���=�* X�܀2�����\Ԛ�����62Ż����θ<:#��Z4��pIߴ����O"7	X���7��ϴY,/�`����?��b���`��W���b+�8!d]?�ш���cO�"����O�^�P|�괙�����Oxq�� ������"d���&I��N«ӊ�k�'����	`��`3�����ote$�Lyx� �HLh���]X�XT������{�z�yB�	��J�&X��c���V2���'�8�=�g=��r�bl~MHV��iI��V��`R�8� R�tO0���_^|G���$��Y3(��H��_�O%%q�T�=,�p�\��^ X�M��崦iM��T	?'i�Ir�
������<��7TM�>�͘�/�#�n�f1�e�(j���9�N�RCv{������( ��_���ӰW[�9�j��[X��������c�l����X5D���KY:g�p}y�	?�H�><U�z-�Ia�c�����p@;Đ��0�C�S��)�8qEv��?���بT��&���~qu���;U�����$�	�qp��K����U�IKK����k�Z�� "##�ml�:��Ͳr��HU
�__R�5!to���~���Qy��
���5SUF�AX�����33����m[�Z�wv�z���g÷�M_����1���1����V�I3qbr����ݕ73lvq1�s�煓����}�X�`�R���l0cA��fi�`(�	��x��}���E��g~D��vP ��w��8�4��E�E#Z9XB�M:"��t��I��T���E-;�e�n���{�m�}����*@?�B����}����>���f�5�PBEwi��(���L�Zj�e��sfc��Nt,[:��W�9Y�v5�����i&�}��o�������w��˔-gy9�G��y��}�|w�%�{?�cʧ�y"�|��_\�����`�Hэ����z�@��>� �^�����$M�&1�L S#��	F��4G>��U!/��"��Տ��ܺ}h&���D��A�քgM[��`�����<Z��������Պ��͡�x!�ϡU��S��������1���/�jFC�F�h�u�dao�RMpn�f0��~9H��l,�C�T��	�z<`_]�(��ꩁ..Ӛ�ja\6q�C��3.F~|du�ӎ�Z��І�o���h��x�.�wȏ7)�v|S�ɷ9TYVT��UTc�e@u���1�3ʧչ�
�T��&�9"��1蝜����^)O׬̭�a�0@9bM[-W � Y�^G}H�\�BD��+H`�;:'����y�[�Pmy���ƞ���՞��6Z�Y.o�[����B�g��x��!�Q!uh��M c߲�.��u�����C.��<�������O��2�o]BY��t}8��m~�שY*į�
�Ӈۡ����r���jrxum��L�1�v�"ϭMG��2�G]Z�֨�K�f�6�z�_���%!;=�y�Ɏ�!&�q@!zx����p���Y]S�����z4���*��3�@%�8v9٦
�&�����Sn�l�{�AR�[2�qFS�S�o�G&��t�x��?����Aq���Dg��B����kcU	!�$����՛FyX��8�y�?Ѳ��>M������l�K�����!`g��,A�?���Q@Z�|pw���Y����\Jk ��<h��́�GԜX�#8��u��?k�Q	5֬ ������q�cd<	 ^W�6-��8�>ԕ��,���F�H�^ ݐD�W>��6�ﭘZg�M�z$T�#�Һ+J��;�̔����ЬE]��]wI���k}��3�_::�eG����J��E��2S���;o˞�4���r�9��	���~N���V�Q��?��ﺝv"�X���>��NH��>t����H8���8��Ǔ/f>�#�ZV�B|�������.|n���&S�b(E3�H����0��R����kncOXn.�R@�i_Do��p�bP/P���r=H��ǋ����i�rť~��϶�;!�ډ���+=�.g}N�ٟ��������^��u۝ɹi�t\P�����~9���pv���:�h�G�%,p�D�1L�E�}�.Y��X���;�f�jun�ʎش+��8��V�`� �m�.N�+ݐ�oݸ(Ҕ��a����=�H��Jm{�h�i���Ū�C�PC�|1�d��'��7A2�D*����0Ojhs��<6��o�ٌ�D�����*����Ca���d����g�.��7�N��l���h:m�.��9d�&~�]w,����W5&�U�����p҇�����E������}=���f���9ݛ��]9�G��F�rb���˃g	��:O*󘠣n��U���M����'�g��y�������,/��$m�'eSB��,��X�W�/�`Ф�ى��>�M�x�>�>ƍ`dG�ͣ��
Z�+�Pn��ܿ)ذ���y�\�|�K�y�.P+p(�P���"��6Ѯ�ѿ�e���k��7�}}�坋U�t��N�-yd��G(y�(r�!�g�?c�f=�G�/�y��%��%���M���p�q��Y��~f�h�+N�2��$[��F�f�V:Iu������@.�.�U뼵���łjS�'��TJ��ܻ�*:c>��~�\S5;~LTA6M��p�r>e���U���VKBs���o$KXr;섔D5���hq.�Ň'���H�따k��>�$�\�����G����%�� >�-��6� �(Ҧ�9{T�R��/�P�Yo�>e$	���P��v�t���Ȏz4P���Z��Vr�b_{�k"1+2�w<刴tJ�X"�C8�y<�<K�Yˈ�{�my�2��
9�D�/��+L�)��OQbع��1�t�Ud�\=u-�O��{i$���Ώ۰0��};�765�~t���.�[�
Z����]A�?IplX����*p]�"�k�<�sպ��Lp��uh�? �D�g;���-H�t�8�/���P�5W����!	#����X��Q���u�P�NO]�~j�!�RͶ���$k���#U�3P���p���$O[���-ذ\jը�7�;��`��)�~�ܨ瑻���!��}����!��5��C�L��s��0bI�>������H+�	`�@_C�����R ��W�5�Դ�sjgJN&�ob=��?�.//���Q�Q]���>�$��U݀��V��u���^��7��o%�I�/.���ŬHL�����������j�4�t[��W�7��o{��j�� }x�i7k�~�v�!y�:��h}�V�.6��`	��A0p�����ף��[�G����O��F���
����7�B���?~PR�J'�Cvp�+y�,��-o�5�+,�����y^}9Y�?�2�e&��O>.##þXe�Ad�1i>��A;����g���3�/���:;WM�,���/Q�.��e�8q���7���AC��[Nu�ĵ��N0΃����j*
��D�l����|�'3خOI3�$�<��[�f�" iM��1���X�6�.ol�q_O�[+,j�CU>+��&P8'�Bvoo/1+RN.�m�q�[}��9���
�^��r���y5��:Z��U�u�^� tPa/ěip|�=�.3k ]�\�Jkh���,�ۊ��u�p8�ǹ����_���Tn�X��qi�d�HM���͛����T��%��P-'��h]��*ˁ��X�=�{��z���5�����!@L�s����Y��U�C�	a�`�RѪ�
�O燷)����OE+���/�#���۞V��F(�B��ada�N�|��	�6'̻Ie5�W�qBN<��;�(�(8���Yu�~S˥,��^�"�}�W�TR�@�
 
�h��s��a;���$�dN����x2q}'�U���β*--���*+ҿ����ݷU��l��D��z�����SP2�LZ(��T�}�.��o/&�(�Iˏ%�{�������Hh�˖d	]����s�;�����m&�Hon	���o�9�=s{Ǽ����I���3�cƎ�$��R;�����q�N¯�	�i�=y�*��#�X]G�y���ZJ�����)T
WB��G *D�b�n02b���3Ч���8�?��/��d���q�+R���n\� K�HQ��η
 �Ub��3�"�!Kߙ��>�4Ϲ�([�c�?�=�AQ'"��ٞ�5n-]ri#�V[��r��ߎ)D��g�Tڮ��P�(�7@�d0fM`�[T�EDuh��� �cd�r��?˔�?;��w�]�+u��̼���4D�@��K�O�8�M'Dr�������ݭӖ�����>��v�#�^}ɥ5c���}����y]C������<�5�K��f���7�te"v)e����Iϩ���KV4������k�M���x#Z ����f1�u����"ȉ2��oG����Д|�?^^HL~%D7����Vĝ2��O�ߴ�Ҍ�Ͱm����p&�=OLė�r��1�o�C���:2��〴���k߱���0����>~���T�UI_@��O��P����c�98��e?��X��^�����£<$@}�3�w�z�xQ4��S��U�-��[^9��|�����u�9t��4��L*#O����b�-&A/��;w����H�����
�Dn���!�H�W�]}|��N�f�"���|����zG��	2-�'v���N���`V~2Yy$�CQSK��,"�0V<U�	�{LBgG?��>��F�I!b&ܻ!��wYc��v��LU������\r��/6X����]b[��Е�{�0J "�KK%dhŰ����b�������b���8E[ؾ�z�����n�GK�ͥ�������݄�@��&���-כ�$�{PK�md�����F�2��7�
�m����H.��x��3;�;�ˡߖO�ش�Y��Hp8�äU	:��1���\��ׯ�*��|���ĬvmG/��K���t]4��0  �gw���tP��\����U-��s{N3�z�w�p+d��(ZOY@�T�`ex+�+)~�i��p~���6���V��"!u����[���B����au�f�z3�50�M��\�%�:�>�n�ϳ7�^�rVW&6���: V���p�^�Qj��w>��ዳ7S�l���1�"������	[-�60f�<��I��Ԣ�n��]V5��z!D�Ŵ.�7}���ZC������5�Y���a��̔.V[Z�,N�@��L}HH}pT�F��r�8���ð������c�A�C�C��@Jd��4k�̾k�a&~�_r��g2�ޚz	�ˋ���J��pb
���#�ا/$EK��(�e(��|����|��O0 ;��Ai5�"
�ĉJ]�)���ZG_�Q,Ur�rK��r��IϷ�D���Y��@���Y��D�8�Y��4n5�n���/	d?\3� C�duA���muU�gѬߺ�,�4�?��~��vM�L����'��z3�m���2;&8U���yz��ޤ�By���Ed7��1�$r�g��ݱc5U[�5�D�N
6��#��ث�Y�Q����v��ICBEy�|����݆k�e/��n�:R#ejO�G���'�%v�?����NV΍������u$2d��z�S�	��_�ji��$�?K}kȴ�o"~��-�c=�E(�B���G},��Vw�ӊc� �NE7�:�G�T�6���K�1�ꠠ��ao��I��n��H6�C����Y���������}�z8=����u��XF����C\�P
\)��~k�>��~�
��*q0O�R�\{rF�Q�-��G�����[.��gve�\��ap�ޮ|5~��o����� �̪ �
�N� �d�~�/�s�w��:ǣ�=�&��'�sZ�U�?���f2w���!���М kmk#��՚).	Ѯ��2Sˬ�P�������?M����5qi���	��f�(������%J�8ϛ�q_.��{��Z�q,"��w�r�\&�8!�8@Z�[%�j���R��������|��c``���k��-��M^FP��[1"P#��
|�;����X�g�	νL�F~0B~��\@18r	 �- m���3L۾��M	g�<����^N��"���l��Kx�kV�p���-��v��J�B',@[�%%F�O��Z�~��h����L�6���}X�b#��p�ʜ~I��M�C�S�KY�i.��	H!�'�.*B���J}�r�{~^�����N�mꃇ�3����K�;�Y���~�e�2�~F�Z'�#�E�؞�� r�A2sɯ蹰X`���h�\UD�Ҋ�-��[}`R%r���]v����M�o��3��Q�Q���X���� kb��+z�2kA6�h�i��^4ێRh�~��`��P�)��C�:ɣ�XЇ�X_�¬]֦d�;_"w��l6
:my�n)j POcȩ�-0�<��kva���J������r�M�9��ߢ���;�4���z��1Ȅ  �!EGT[V \�2F�r�"m�"-�Tl6-��[z|4TTT�Ӿ���N�;�T,VM-����� ��K���cϑ��6��&[$ٚ��I�1	�����T�}��+)�aav�͊���� k�L'`��s�ʟ��X�txMGI-�0���K^��k��C�b �ߎ�5]�C�;���uL��+�F�����d��{ι��:���ou��U�L#
:�����?��G,&���8����m�O��2|ݾ���^Đ���B�a9{�y6�K�`gU�6�����x_�Z�OUMLH����n�԰?�qF��f8�Rd'R�:}F�h�>��fͦ%�L�Az�%k	*/�Q�xXw�b��&�#0� ���.�.L`�|�^��χX,-�~,��ܷWVߓ��YVP=[A"�L��a�Ep����&�vla�)���I��d�,FR �!�&��\ɪ��w��#��cᥫo�l�|9�m���(�I�8�W$V|�d:\#���Yv�}ĕ��(!$�݆��Ƙ�633�?2"���,��M���/>[_S�ۖ�P=ڂյ�LFF�۽���%/�.����n��x|~=
���E����%���|���}_{Y�Y3hJX���G����L���S�۞4%sae܇��O��{q� �~�J�To�a�w}�rĊ��?����T��Q�S6]9m#��{���w%�B�c�dW4�.�M�Ԥ�=:$:W/�`I�9b��U� ��n�9�gP�= \�J[���ĭ^����h��� �x��I�y$]u�~Ȓ�^��v�����z�2R�rkT�y`x
{|oϷ}	�@�����h?~��?k��F�_X�����j�^;.!�Uß���!::���wt�gnJ��WY�c7цAi�@�lF�Nx���29$H�#�"��"�**�7b�՞۞��� W�1��:[��ǡ�]ă+KϢ^^���.[{�?OF<�$���Α5 �����T�֙l��+�wD�DZ��~pm�8P���V�M��`x�H;��k�F�sO3No�:F�!�Y�H7mR��6�}�5�KȦ��]�(4f��;W)�JĹ�N�������ί2�HΌM��S�g�9Rnŋ ��X���5��pL���V��|`w��e���`��Pǡ���3�&����:�VS�zY��z/�9bUE?TT\&a���c#<BB��� s���q!}JGU�����Z�:�d,|�P���T�}8����}����'y�)��)W��V�D� $��jRZ����y�4��&}7y�D�∧4�5s�ab��L�7��s������M4+�4_"�����Ai��L/~��߳탏�^��#��p �"0uCW�1�l�3�0����>�D_5�V�ww����c�9�I"�/⼁X�-T�X]���T�Q�/pƁ~��0��kF:�&�r8�ŢBf�ص��旳�X���5Ng�)��uLku���?��O�C�f�,��u�F��@4��k�?'���$�<KJ��}�,�Kwv����ǰ\sS�Hq�Z\acVnnnE^��D� ��ʡ?�+�T-jŌ����g\�$G����t����v�n�3jj�cC"2h�(�󹴔kׅ�j޹|�
	�n]�{=*<K��3��Z�]��&B�)��l[|��.c�o4X7vz��8�����ᐸ���(�KE�����Վ�޷+?!UN�e�Ybԁ�c�aS����_���.|�Q�$A"�&D�j��nZ@7��M%����b���k�9���>j���'�F`��4(�4��|�be������	%�D�P��������.�J4�j�S���|���*�S�r�%�❖�+Uԭ�0��2�b#$"Gr��µg����8Js������Ș4��KW�up2���w,��$��%�k��]�Ω+�����Q�<���K��pk"��䣏?;?� �T&��4��@�'�����+�Ե\��O�������ſ
U�G�	*֯���N�����mh'��`_�^:m�Z�*�)��%�tΈ> \!��6�ζ�M�`��� G����
�>�((?[�.|�.��.�c��;_8�0�V6�4!V)���N����S���nN��[��ʁw���}�y���s������1�K�?����`u�o�6=m� ���B�_K����݆՝`���TM%�P�;$^s�՝��l�U�|�[�[ŎB�Gi���s'���u����k�����<b:\��`��C�fK
�SD���(�-�+#�n��}�RO:��~��|+��,z�f�Wa��)ʪ��,�?�
K�u���2��_E��1ܹ�����������H�TD�X���[	}Hā&�C���t9�v��Ll�� AH���gs7g�����\Ǭ+~
N;l�'���w�5��Ė�mI�����o��A;�>�w�S���_��@�O\/�A��W�v!Br@���b!�����}��650���� �6A^`�A����UPitK`(���p%�'��!VTC0	�G�m�f*��m}�9����\�����ϼ ����������ϩ����u��I�9�o�x�����c�;o�������K�>�&>.�]�+��	�^�[��6ܸ�e�ή�Ô�j����#� q>�sT��#
h�� |'���,�ђ�!J��)�Ӕ�U<\A���e��ȗ���k�F�w��-Ƕ��Y)y�w�]�u�ka��'�I�u�xz%|zյ��N�7*&�Qu:`�83���N��Y6b+��z:kM̾��j��e���	�s�ٳt����p)!ae�rm}w��9N������U���z
b{�TEt/g�xw�p�vO}d;��Fٗ�Y�o�UtK��k�G[�\�C���f��32���<����y��\��`H8���b�h���M��N>����x]��A�Jh~u_Sj�]�&����'�^��GS�[s3ف�=��戚�B�ݒ�;��&�s����p*�N�������2/1 ��۟��Y����>+K� �	�]������<-��|X��I!J�r�A��F#	��'t~^'xL��uY�z��'����Ct/�F�NVW���_�9���V{����_zW�)�	��ȷNf���/�o�E��G�^�����#[��o폡�;Fq�k�']�徲K�Ĥ��`��:at��$L�}c�(3n|�W=�up��~n��ym�;���$�����='hK��}�-�����|��N���F� �� ^^��9�������+]�қ�ώMoBr_��c�M_,o�pjK���o���@D���@�8B�88�ɧ$��.z���c��9�48�8oK��N�y�}��{�^�z濰��l�׹�ǁR�2vO���_VE�U���lK�OX]�7�K[]�Nq�����\�O�cl��%\�S>����������Ԁ$ۧ�c"k�MM%���63��
��L�֜��U	���,���t�gC4艓��x���K;�L�ꆂ~#ܹ4�c�-�n�f��H^��4��W+��'f�Y�Q��qD���Y����=�����c��ΎO�f��?_G?��|��+?|������ŋ �!��K����[�eѪ���'���ڽY���m}P�<�/�}�"V&�����î�'S�M�2���,��F���":�~�MR��c�1�b�c��'��3�5��G$E��H�w'�Z�g�n�$��^�U/����ꛑ`�\}��9�o�߱��*�|���?��
�/�:�QALD;�� ����T�y�h��j����㺆c#��;l��LaN��K%f'�3��<rV���g�@�-cu/2tC���z�'��y$}T	Y�8)͞G��#�;E�K�-���;n"gT��gS�l�v)�iƁ�~������<bl=���������^���� ߰ �����n뮃c��v�n��U+�`��w���� ��5D�Rn4L]Gt�J������>j�C:
�~55x���<��0����,�af�PVQ�4�*v�P��H<6��pE>�_��]�",������ko-PmR+��,�T�4�L�}�?�\8{�s��I������r��Ov�cGV�W�c�;4���	n9mD\+B0��`+<"���`���2����V��*���!0WR��5\Rs�.SICVnOq�c�qi���\4Uev�y��!lȈ�FL�l��	��L�1}Z�7`cѠ��Ia�;u���u%�� =�H:�Ev�8��Ov&*���j������bK[�����LT~�-�=����0Y�p}��d/�.��6����t�N�NB�mm�V:���<F5���㋑号�7Eۂ�����l�c��o������#kHZ�Å��ed���~r_B�׳����;�������-�P�IY%0Ґ`���C�<i�J�cEM��a�:�W�^�/@o��}�.�#A�V��H��_Ϧ@�|5���T�����f������Er*(m����-L�_Ɯ���bZe{+w���,�p����O�������UU7jJ���{Ο�'���*Z�9b
���	�}3{t�}�T�~4��Áh�s���/�;��ٴ8�c��kB|��G�V�r�vIl=%5Wa��E #<��� ��X�{2�:�i�̡��Y��P�r�h����S�aD�/:�gc�J�Dz@�����Is&`=X�S��̛�4[1��90��gqmC[���z`,8�S�k2N�ی�* ���0��9�"�Za��Vì��	�0A3�iX���������+ض5h��������Kpwwn��,��{pw����5��{�ۣ��ڵk�Z�U�|��=��Tfٹ�Z&
�𻍌"ʯ���`E
��rL&��>K����䑂[b����|%�Z6[��<^_�:��M��"�~��:_b�7��C���r�����h��(�4�ϧ12���Ƨ 2*��~}$�9��st��XPhU{��-���g���d�ni����,2�����S�]=_��p(m��}������@��Ŷ"�h|AB(^����gr�#M�3��5 M��%�����a�v�Wx�=b��wc�����1������*
���g'?������֌LQ؍W�Y:���~^#��;8u$.(`r�P@1P��S�=�ͨ�y
��9��)����Yw�Ì���X �����%�i��3Q ���P1h�����[�(�n�O�|z�8��JЈ@mK7~��������!i��$T ��0	��Q��i!0� 5W�\<i.��I���'6��� ~��Ч��aE�	4i�A��7B��`����9��������	a��68 W�D8T)P=e�夆�oݩ��cU�|_���~ 6���IB��������G��0����nr}���|f&dB��Bٳ=&=-��c�.��a�D�/BA��ŠyshJ]tWV�#�Qf-=xO>�J�B�{j�Q#�;|-DI��!�����-tȣ����G� 0�7�O4��H�Ͽ����3��D�a�x�[�7����݃����W#d|;mh�;_��u�w�\ M���=�[2�hC5����p�l��Q7n���\�]� �L`�lȺ�toH0cl����Ǘ	�A)	�7�4]$0l���8�_���s�h��]K���q�P�nKE��ۮ���;���|20����M5�p���(��翕-~V���v"��3j<�f���eC�B���]l��֎n	�F0_��2c��& )�����Vp�ZB�4����W���LA��nU��_�~�����>���;�}W�ȳ9���8ކ�m��ND�U�ז�/�<�y�����[�=�<)��v���W y|������:T ���w�^��[G>�!Ӊ��9Z�j-s�'?�E�p��0<L�^)�8��?wU����0��5e��;ܾok��_�*���\E��ם��ʵxl��M>�?v���B�z�a��>�;!�?Ў��s&�]U�}�_�tB���8���2x����s���i3T�Z�S�W��3--ٙ�X��]�<@B�YW��6��C�<p��h:���1����cպ��$�|�{���F\h�o}�w��a���Mڦ}3��������싢/��}���0��BЕ�]�Up/�r����x���?6M���8��	r��	xx�.Y�2�B�f�(�}��-k��6[�+Ǎ�h9��68�̒�(�,���=QE{�����E�Q�6����y惝�d;�HZ�P.���޾���1�&�u��0�L�S�^��M�/2')��z��W���w~���n�&��z��*��P?�����G�HS21,�~�aC2VW�х�9Rb�a��	·7�؋B$�L��Xm<t�Ž��%�/Gkq�8VP���ݠb�z����8S������E�)�?m~�Wq��U�����>�G���$C��ڼ��������{��W4?����zSo-*�Ƣ'�_���yy���9/9���ͱ��8Κ/Ֆ�����M�l
|���Ю��]E� �¥2�|��"*I�d��nc ��P��O` [R�|�)-�`���w��Y8��+)�_�gL6itt�rc`�M|�����A�(�<.�;D�R?��=/��ۙ�-R쾗��'I�ĕ��������ɧ��l����s]�M�Af�}�U�ǝ�n$��*��Ҡ�N,��)��`����X��[�8��*o,g,���u�[YL.�mZ}��캓Z$o�a.~;]_N���i[68���/������������Յ?x�q�~G�o��6��ﮥ�V�~#o�_pv�Tgf�ǿ CB�\˃����t[�b������_��-���|���%�lx�7$�c�Dڹ9��&�:�|`k����g&��1�ٍ�Ec��Gs�����ꓶ���:̺��JA�H��>41G���p��RA7�5:��{�u��`y0��f�����^����	���b�����0�ĳŮcȕaĂm�
��2��3M�H�݇���:��FZ�¢�r�\�1����=1�G��0�����̾�O�s�kSQ�x����5���I�ϧB��!�����<�n�d��g���Z��`b��3}���)_�����@E��/؞�\��18.'��#!������ֆT���-�� 8��%(h+�y��:�}^M1?���[�^�%s�d"�D��c�%�=��c���=�L�l��'�
��f���W�z��M:j3Pa=�i�f�1�yo�@m�c���2-_Ӌ�^���x1FM/�j����Hpjo?q[���з)A�xի��?��S�����h�ŗq���{���K�ٸ��Γ��>1$䅶.xf3�3�[��C�kKۃ��`#\��9���NS�N�3E^$���UPж<=޺p�Q�F���n��M�]���فr�Q���r	�.��Y����b��L��9���%y�@N:UO�g�;�A����yl���8EC�l�<5��CT�,/�ܠ]��2Ѣ�S2�q��8~�3`��I8�����O0)�q�LNK��۸������$ݦhoo����n-�Ϥ�U���%�x��H��^N2�M�,#����=b!��R�H�c����g���S��Ί���S���`��7!�����L&�s�7��.�Y6&�f��rd���p����B�>f���6����i[MF�ЪJn��=�1w��oM����'2���7���淋�!��2G3GE���������f׳'��_[yB��ZE���	 ���"��3>B0�^�_�.��v�?0fX�� ]x�D��~c�t�i\�@�â�jZK�`������e�]d?���w�uCկ����aO�-%����hdæ~_u��'�պ�BlЬ�8�WU|�m�����O
"���{�q7Z�T&��-��v*A���ڸl��}����΢�|�������7Uº%����A��,�o��ژ6�I�aH/�A��	��_����΢�Z�7����=,�����$Q����C3h6��a���a����f��B��Q;�Z6��[�&f������HtV�XiW=<�s�\KЙ��{Nr��	��X8?�--����}<�Wzc5�le��^�o�x��DL����Z�Ԝ��f2��$��T��\��^G�<��HS�k���J��������=0iɂ�x~����%�΂����z�C53=��W귎����Z���<�lx���Ϥ7�S����M����U[r:X�@�ruLEc��ǧd���A���hPS�6_8�T:BB���5(1��^D�W��X¤,c�~�n��B3��wg�<�H�յٳ.Aw;����>~�Ǔ�P����n�ZO����8�w}��y��]xt:{0����#�߯�l4�=/���'���ss�=t��N�>?��[g�QW��)����ds�D߿bC�h�A���R;;I=������"�v��q�_����!)�E�d�����K��)���r��^�g�c�軤V
1M������`��w ?2V����wZ)��5O%�	_��t@4���������}c[YM����\�m֛��<y�[��HwP�R���)5�q����D+�}�0q�m�|����Pb����{��͞r�z[��y0��}x:&A��ġ�ϧ�еaӛ\�!R��A������IXCpy�����Ug�:2������^v���S*jg�>����UT6��s��V?k'[�\/��H�(Z�����pڼ4�r�qJg�9m�Yk̐g�Oߡ���:,��G�EɾS�>ܴ�["�ם�@�<aO=z���L��\Y�f�:�C�pm����A=ߜ��*��P#�2�2`�k>D���܉���Pf�me���w�1����uDXX��G��BUS�ϫ�0���Qcp5D&����B?u�k\�2�z��F����*)�a�(R��)�����������pY���G"�jȅ�'v�C��	�̥���WDS���-|\����;Q���ʌ�g�.R6�[��}�}ƺ��Ѥ?�K��n�J�W�'�)3q+�W'`A�� ��vv��P�Dv��bg 5�lx���������i����͚�������63$`��F�7��X Z�^ߘ�cc=��|)����� ��4���BD��~�]��	�ņU�25�O멦�o5c����a��R��0hU����Y�6��Qf}y�\oN�R�Ȃ����61��eT�շDL����_�+p;=0U�)��8;UxP���#��ϟ�A�;P`G�Yam߶���e);���r�}���!&p�O��%���tӿ����ի��rc�#U�Z�;F�pP� )~�����Zs�zI#f��^��h�������J~���C���F,] ���w�'%t�*�W��^��	v�YFaG��N1]���}P��Vb^+ԏ��0O�$A��J�������}/���p��/ǅհQOU��i����T��:�.sDĠڳ�$�}�'����5ko
P��}:���$e��_��CC���g�D0�|�@?� .!lbm�ձ�e�k�}��٣����ބ��������ᶜ`�Y��AY� r�o�
#�f�<H�CA�<v'ͫw;��#� */W�e�����+*�sCo!�ǥ��KC]�r�ȑ=
cAB8"ʄ]��p��7c�/f�?�Nѱ �E�{���l�4T�Sn7^վXό3��9u��3t�͐B?_��)k����W{�,ڊ�@m_H�W��YLb�w]c�V>FX��7��8F��7������H�S���7���C���q�"��g�:m���M��C;�_���P��mr��1�Z��J%,��9ズ�QOV����{� ����;qm9O4�i���I:� +&Z�]`d���M9�' �����L�u��߹��82o���ݖ9REn=S�GA��F�)�+���X��2�[��\��	[�"��5�}]�=�VZ��@���~��i�v�<Y��}�����N�N6������E�V��P��lU�"*Ԡ�xW?zσ���W���. �`E����C��}>Uάԥh���p�9�'���,?�7���b�0���D�mi~�S��۱�"AK�ڬ����N�o����+��p�lG�E>�^�,�1��+�����2��^��i#Dm�k��̔:��t ��;�3G�!딲xt9�݁���.�Ai~/���3a�m0t�+�W)�f-?XR�6��x;�?6��	�� ]I�$1Ƥ�"�䱟�mA�ZFf������+PTL�e����(BsNC힉�(��!5�]&�I�%��+j�+��>{��o�V�a�ӫ	B~d�~��ŭb�D��g���s�]^�;�_1�����~:��;��4�&c�L�Gc�7�w���9,�o�"�e�!
fbj�Jk��S$�0'��kO�Ō�\���m��te���,rm�"�)'����	�V���G�iA�����M�R��1��#���&��8�s�ؾh2�E��c���͏��A���A��E�T��Yk�4qGQ0ۺ=�sv�N�?��ǓfC��tm/%��q���{����s��W�gJ�=`,��t��v������~�)>�e˗��.Į��XM��e���P���z��ڄ��^��������$�����Q��a�*�KTѼ��O�+���G�h��
m��L3^����A�?�:��6�������U��0����x-�:�����m�9�������/9���	������D��u&���R�}�� K��l�v�z{�+ӎ�������v�;�e�Ri�M�rfx<T M����tT���+_�}�"��F�>���Wm��6;�g��8׻=�d�އ�E`eztˮ}#�B����f���P ��{�i�蚀zv�Y���"�:�����~�k��Hu�}6|�ʋ��aj$F��w��|KX�H��ن��@�3������j��`Ɩ�sB?�_߈�
���B8|
���IǏ�� ��R�y�:LgOC] �B'E�#k���Q�����w�د��	�}�n��}�Jga'�Ds������)�U/9"f6�[,|�Y��~[��hWqT������ �ˌqr9Jʤ!�
����m�7���i-��]�A0 ���Pp�M��;R7�(�	pbR\��g��g����R��6�L��Ի�N1G�I�G�Y��z�oQ,�p~G�Ξ;�:�S��#|Α�X�8o�g�U����YP��hy��3W���A�\�x����ʧ�r���:�e��w���7b��r���PP��inN�|�ȷ� �ԥ�i���:��"�w��Q�;�)߫)i4a d�}�Hx���LQd8�h2���|�u����oL���D�*9Զ�"*��!R�h�C��k�a:no��sB��S:��b>�^�Y�G��4��`����n����{Em,���T�$Y��WBպ���}9�X����?�i2�U��BD�aֳ�������-aG�=$G7�{���=(�WV
=�wP��L.�na�b]�ȡV�*����~���
�[��e�����W3(E_��/�݆�״�N��2>ګ�$1�)>�E'�惔;q�9;�c�,mc䵴���`�+�[�]�F�����D�Cp��z^@?j��s�RN�5��4m�Ӥ��9����u��^ǲ}�U�gT�fk?��{��;��I��9�P���v�z�Mc�4%���=d��0��e���Z�)Q堹t}Z���N�W��臢1�X꒿�e�)��5o�I��^��1���1��D+�l�'��s�YQ3'�z��CBd��G?�*m�Z~�~��K���kG�=���Lw������3̊��.���w��ٝV�^CT&;X�-a4���F���-j)54�T?Mk:��+^�n0�m̘G��e~0.�-����RYPW�^2�� xO����@kX��(FZ��d�5���/Pz~&�S:<���.|�h�l��5��t��U�aͺ	j��B�wͼ�}l>#m�������Ё�d�[�-e����%�r��/!��v�C�ߙH�h'
n@�wo��'x�^ାv0X��'���&���7��|�z�v��{3��V��cq2hQ�<D��ypq���sL�,��C��+��Π�J��&�K��*�]1Nt�i��0�����N�w��N�r�`T����{��)��1^F�-�j-�F-�V3G��D�~�JFp���6z�O���D�Vjxw%,؆5�g4P"u1l�e_$8�#���~�&���wXsBw<��>�V�jM��!@�Ce��e��*��9�N��sXfȲ��yȀ��B�;%�O.!L^�=2F�R���8���"tUK��x��a<dy��f�.3��[�嫉��:�") :ER��v(M�k\�;נ! 	y�4eϙ��z{���[�h�Juj�ڷ���`�n�B��Ⱦ�Ц5��2 �����l襎&���2"�E�k�:/�J�����=�6H�DP�1�i��T�]6Sǭ���o^������ck��99N�K�.��]�c.eh���7�ض�˒Q?��b��׎*�[�X�v0b�~�ԃA���6yh��~�x����|`��H�B���q���U%W-��3)�߬��H�o�J'�!�E5q��x���m��ߦ;��^�F�����N����\�b�O���Q�z��ї0���r�D{箕��Ҵ?����Ya� x)���8���m��~�7Sr�&��"([���C��rqa���f���I��O
�K�"Ơ���+��P�_D�p�)�y2��_�-ޘ��*��nB�!��d0��/,o�>�5�am�{�D�6�5
[\����G�i'���#"��]���m�״*4�������Eɩ#!�g���88�/���Ȩi����E���;Җ��w��@�0�N�=T�9�B�7L7@Qh�{E,��B�	���JIG�n!�x�N��f�*t�*t�ز�)d\�\�1`�J�$`��u�S�r�3�B0[~�nY��iK*��<��p�0u-o��{,O�P'�7�#J4����O�&�;^n&�v��_���<=g&�L��¥cs������I���q�x�Q�_�.H讎3
��L,"{���@1=ɓF5�pzd�>><c��s����A�?᥏�6O)Я��A��%j��Q�M��G^?���7/�����o����`�����p��.^�=�TY�g�x��D��XT�
(�	���� $��D:������M&��"_����%l�sP�K�)\���p��G�����c15(�A]�*�bi��-��d��R����'հ4�'�4��@`<ko��jO�PI)�W�J���^�8&�]�k5�p��Z$1��o4�	�	�X��4p6�A�:�*I����k��G��^�e>b��c�/$�d$+n��g=��(I�I=D/��Y��u�)A}�9��D�<��e��eIۊ]�~�g}h�c20��?b�IyEE��q��O�_x�Ya���@E(1�+ �f81�޴B�^�B#�ی+S�W��5��aZ2T��]Mik+���@Iee������]�w*<Ol�ȏ�iC�ݼ%S�F�[����:M���f*I=��"Bw�L*X^p�;ߑ����)��m`��5I�rZ���*8�yGc�%5�kc9���
yk�x�_��ߋ�'u��ª�i�Iv��S琔B��G������D)��l4�B��8�8�w��:���K��:���f��^�S-�079�:�_��+D��+�4zL���⡗'ü~�w.c���z%v�+�݋�����B�rV}1��T_�S�_1�[5���c���;p��*��+���2� _����ݾ�U;��c?�Ca/]�w\�K�ʛ<F�AG�`L��6@��ec+�OTF >�6ҳ��+Ҫ�����$-s�����g-�p�=k���`��K���L0x8�/\r�������`����Ĕ�LїI]ت*��u; $�8�b� 1��0�Ya@)5���H�<��% B���\(�D`>�o�4�nfhH�g�l�]!�r�I�I�3s��g����ڳ��;!�rܫ91u���S��q����hg�DAs3���Y��1Pp�bpO�MKKIi�cK��f�R�k^ee���Nt �Ox���,<�sf�:�s�9u/��#&p7����P�����#��f8��qK4��%�����<,d{���=C����Q,g�=�$8��d.�ç\�
V�U��BbIT7B��Z2�V�����E\�Q(]���A
3�&�C�Y��/������si��:'��^}��~4�-�����,8�R6<�&4�@�A�;K����6(o�M�$Q����1�	��.^@x���zN�n���*zv˿�>=����욼|�Co�>��M�/f�pCQ��gL�秚�+W�d�,���x�i���W�IN�B��z��'�˒�޷��K޺*#4V����(u���X�3�P�f�9D���:��;::_ltLwx��q�����&"2R�Ņ}gg��Y|�ه�uT333(88�E�4�����y�B��X�37����#��sVߤŝ�PUx)!�8��N7� �Ɂ�n��f�AO@P�h���Ҕ)�7_�9K���<\M�����yNU,d��\���s�?���N��o���i}���͂�JԆ�!���=���4|�H��á7�{:&8�>fy�eZ�1Hi��f��
0K��b~�F���[U#z�^h��>����x���T��kG��c[1'I�D@���}�7(U�m%�� ;�Ǥh�2P%,W��j+�ڣ� 2�ۣ1�'�c�_�{��7��bP�hD�l��M��}�xw~Yۣ�`���^J<���;�X��:VD�O�{EZ�=E��T������fJT�a���:��g1(Pک��d�!��v�6=�o/꼟:+�:DnRk�$�ݶ�Z�/{r5o�~�v���K+ �+�W#�+�Y�m�gi>Y#�jiU�*�{7Wό��ᙘ�W`W�p��M�VU�⍛,��n诮%ڢ)#�p��������>���8'�t�`�a`���I������B~5F�NJe^ѐi�l%ā��7��9kI_&o8���q��O	Қ�Z�x�@�:[���q��m��y��y����d2Pah�8v�P]֡��l��Ԇ�p�!'S��Ah��C�>7���G�dce��8Ģ�I�}�u�C�ǅ��c�?m�_&���\�������)E�KKJ3.bz��}��b}��sV{N/)F��0���>L��+w��h�N�Q�_�/���&�N�yh,u���ϋ'�B35��[���p�s�F��L�MMS�&�	�$u�+..\�|�@PP������@R��T	*�=��ĭ7�~�8Q��ۿ_z�5b��~7G�����ݫ���ၰ�;ZZAƆ9�'V�N�02�W52����ۛ���*�)S��V,��i���!p���Dƪ�+\Ƙ*e�E�^T�E_�}&����<R�?h��n�_<o�K����/~�vU�()�d��//��->�+)�O\=]�Ƚ�C�{:Ė��;�[�_���ū����������@�/7/P@�צ��dP��0ՕD�~�E>��l7o(�r|�=�ٔ�ݒ�.Z���:7�A�;���᭷�S��$��՞��@kv��a�1ƒ�F�|�t�4���t�1ޯg^��[>e��� BS������É�?�M�V�w?̈�.�z3`�[֡&�R�g'����>�\�vY�r5}X��ZN��qq�P1i��k��|/I��k��M���O	�'x�"�X7�_��3�B�sQڅ��n#eE��Z���ux]Y��C����zg�<*����-���mAB�������i��D?{������<�l��쁋�|�g�������~��=��2���	ۡ��%pZ�8����]�wL�l_�H='������ڼ�z���:r�EP��mf�[Q�i9^�R�~��k��VVsM� ����a��N� 8G��$�p�.PԺ�y��:=fa���r��}���4ZZ��,�P�b��Y/D���K����^��"KrrrbFF���'n�{�13�׷7�a�S�f,W�x~�VC;���f������Q������e��esee埻TuS,��츈NNNJ�NS �.�"`Ǽ�/�~� ���ӎ_�b���ՙȬF�\qyƎ�{����:k�%���_]pؕ/:7�kUG�JJBo��ؖ��ж����%n�x���W;_=��j�>@4~{��N�\�rl�R�P/ ��E�����ە���I�H驣Ä��n��k��#��P�D�7Y��m��=�&f�7Z�n!�.��@��h1����a�+]�7�� C5��	s>�2��oa�W�DB�~0��(uR���hE���p��*Q��Z��u��h_��o�M�ݩF�r�(����5�}�r�G�蟁�����G�2kџ�1ZB�'.iM��\M+�C\|=Qe~�:P���x���o����WW�[+�w���"��iF�.z�~�DI����{�� I�������*�.X,� Vk��E����8��0M�c����Qu3-醛(D��.{�����c���?|#���y{yx(u��N$���.MBK��H'G_ /��i׼:*�(V�Z�KD���N1��ҒFZ:"x�x`Du�ۑu�b7s�;m����k,���)�͑�lY�ҷ�}~j�3���\\FB��w*��O�!�1�6�(��V8?�/BT�?ܣC��Z<ܯ����OvC���U9_F7ԎO�O��/���=O���rQ[�5�Ɠ{�~�6c��gGg##���|�%����Æ�Q��|���W,��3�=�'0��`��+�݇��lf����^7p���_s)ɻ�{�	��:��6ysנE�H~vڞvz��C���z���H�Cd�j>�u#�W_cUUn#N���DcM�س����j�~m�s�.�1�n�3��q���t@V1��l�Q�׌�3��+�����3��5��Z�5lY�P�79V��I���)UƋ�:�c�yAқm���ҪUk���v�W�Dhj~|&����76�ѧl���$t�J�X���ٺ1c�G�0��o�|!d$'V�y�l�"��be�ѬE��zmn�
���aF�3,�--��-W�.�O`��;���dw�:�{��=#��6� ��)vn�g��[b ��fUkkk����H�<dh�e��@�j�BD���E��B��n���>��{o�#j5��dB��2����mV��6�qؽ��ŭ^�ԙ��2p�j���-�:w��J�[�kTZ\O�P�4�~���e1]���$���Vl_4�`�F�]���IZ]���f/�ZJ���D%�hwI[�ԙ�U�Wx�v�@O0+M��~�^�2�@}�ӏ��=���o72������!uV��@,�l���=�a$_�:�+�������:;͠�Q�c����楷/�0�{�Ђq �5��˨sfpPP|z��Ztyc#漺�ݝ��'--n42aȴ���(?��T��.KJ �rp�{�Gռo�K��<��X�����J�ǫ� ����C�V���5Vӡ����#������+6�vP0�l *�������z�ݾ�RE�4��8+j8$
1a�g���ɲP*�;״�}���7�9F�[���oاz���j~����ݽ��ڡ��9?0k�Ȁ�m�M���L��y����f�!	�+�Z���f5��&'��{��3g��� �(؜��o�]�T�2��x<�q/��\t��I���[Ztr��V*�����ф^N*��<�V��������q��Z�w��m�,*Лvt%!i�}ʼ?��)b�l��9���>�c�
 65�NGKG��� iw)��8����}��(��>g�q|��ޏ��E0*�+�\YY�T�5q�^�u��dr`-\�������P�R������|���%XH��64?�F��d��y�U�͇7@vFN��N�Kﯙg�Dݺ�05j�Ə-av�L��1f\�8�17^rZmF-Ͻ���G��M��� .׆pM��U�fb���; ��2
��PVXe.��N��_���fͨ�c�n�Qn�����dX�(�'����tDC��tS̍�V�@
�N��$��\!j-��~#�m�ԇ��_*=։�qe��}�v����Ge�;}m:Rڽ\�'k�.���������ZQ{Y������O�r3al��ę%xP?�" J��S����ͷ����X��$Ә��V_s[��5�nU��DРz-q��s���C%��N8�_�,�s�DBw����	8$�q�7����7�c�W�`^��5��Ut��}���[os�/Q��T�������?]A� k��ף�Ke?ߡ�9�Y����S:Fs~��~Q�������_�1AXT���U�塟��ͅ�Q0N�uj�v\:5�怌�Ah�d�� n(��'�/PhW����B^I�ߞ�%��.�2^���-�C񅏉D�#B�0 ��/~�:���L'�&�fHj}�,�2����@�S���/ɉ�L�U��\mn^��@$�\:H8@f\g�DM�H�ݷ��;���.���ך~�nVA4�xЈ���E��*�V�`�ˋ�H!�|�N�R����ޠ x�C������o�)��lot���~�3�|v�(F(�ܱ��u���o����:,3��OJ�N�m/�!�WUSp	������']����Y�� ����+j@�����i���o~C�4�`�����.��ｽ��M�Z�wp����(�u)'5��t�<��_���``G]�.wVײ�"�Jb{�Gi��L�艕�^��W�^t�J��S��PG�%�Su�c��B8�#ЭV{�/P	��UdC�$��g�o:]�%&����冀Wp�����C�������3���C�
Ç_&��r*~�2��#��ݭ���\�W*=m�R�⠟�
0��&/p~����m���H�3��I0��^8Ⱦ��/ϩX�H�u�����e㮀����h��_�lh9�X����.�L�|��V�[iB���3�Dvٕ��Ձ-'�7c/�r�j��U�r��u��qr�p7�p�R��Dk^��ҦU�h[�4_|.Q(``5�V����@���N�,�9؂=���������m�|�40sp�R�:��7[��.��r��;��9��ҁxź��<�#�|.�!�wX���7*U��4��K�_�unT��c0:.��-� �������a��jiiIMG<�Ct1zb�ƚA�[��&�� ����F�e�49J��N����U�Yv�H��p�CGj�iz*����N� JҦɮ-���m?�b��ΪBoH�<-N젥rY��b��n8������e5KsǇCU%�E���+��h��s���$��p	R��t8��*���W�̄iP52��zzsxD��+�C>�JA�8��#�u�:��y�e�d��U���vf7�Μ+��.��$F�M޶����&]�썹��7\���lp0�B�/+�;�%w�p�������&�Q_t{��q���Ѝe���}��ÀiĀh�����q�E�w��P���Ȕ]-�w,����q����@��W�~o݄��G^1�,���Gm��vx�&oi>�{���+����&�̿&s3�����y���:ٞY�db��8��q��9BH�4�\d����ɶ8��J�� b Hr���1ϳ̇����$3:�S2@�r{='>�>�z �[%3��qt��sMr
"��N��������t�J����[H�9��pH�����M����`+�\���4p���1_4�}ǭ��
q��BU��>��
u>�JuJP$�*��.��;����ZjU��N �����Nє��r=�kÕ6��n׊r
�F�fZ�r�nTv'\r�k=#Y��� ������F�}6��=�`"���b�~��:e�+a9�{FX�}v���������&��������凑�mD��a�#���C�vF�ѦI�uo�7��>�'����r�C�xa��v�!�.�ۀGW	�,�۫�|�ʥB �v��U��J$�7_�6����w�U:$u9j��"��jʣ�3�q~:h�{ט6er�U����Fh+]Ƨ������������ �V:N02aqWio>�ܰf�k�?2)�k�[�:��	�{�31w�ݛ�s�<hs�!"�����&�5��6���A�2)��a�A��}c���u�W�5��VP��bѐ�,�s����#8����q�U���f]&�<^.��6��p>�������]��]�'�Ҙ�Q-�w�>>���*T�����C/���_Fތ��$����WN����{��K@k� ��i[�c��ica�		7B����O���K6�b�nvT.���H^_W&�y@���2u�r����D�z���F�ߓX^%�(xB|����r��b]հJ�:�gOF�H�#
v�~i�(�����J̈sĉ<�<��HT����u�sw�`��!�Z���S!�텺���aᏖ5��T,��@�#�wC�$��͸��^�����>쀀v|�v�ru�L�
���?ؤ>��V�O����1��r�{�%Ϳ���Y;�V���\~��6����a��G�b�ً{ä�LXU�P���b�:A���-�h�gp��4�Y�MN�
?�"|����#���h��-"���Qf�)ڕ���u�;��׀�1�>���o=7���oR[��d�V�`��{kl ��<&o�F#B���o�o�9��Z/C�ʤn�p'ӒT����2�[���*�X�X�s:�oiA-E���l�F%]��"G�AY��r���E�v��S\�!�P�{�*�̯�͟�Bi?��|Bt���t�Е
���@�7�r��mNA t�ףՐd�D�V��޺���Q��}F'\|������'P�aVE�x�c�K��L	f�7g%U2�+�T�6��9LC'�b�~oDs�h�`Ft;&_N����䎑#neE��k��PӨ��G( �Q�u�Jd�)��0����+d�k�� ���@B�[�TF���S����)�h\���������Qc6�۶m۶�ƍ�4ilۍm���|'����{���2���s�^{�s��qЕ�n���2 ��%H����yu��%����!���2��b���#�g��[�R����QV�-�W}t�nU8:�����&�{{ϱ3u�9��Z�����Uh���. &��kN�*�?�����x�"�	�k�ʽzl���|S�̿�׻ޑ�:{�Q��k_5�6�g��'�2������>�� ���$}�{��ͻ�"ir������S������;^�2��kg{E������ԋj}M3�튮�+��%��T�6�0�H7ᵁ�x}A8��K�f��a��K`�!�]�.25D6����W.Cr9�S��ܨ�ᐽ�6s�u{��b��7id>�͠������݊�XM�Y3X�ǧ����C!)�3�鋆����2�����X�+!�3�ȍ��a���p*H&�ǌ6M
 g�F�;���N\�����Ӱo���u���� ؂tuR0�0���<�{X��H�A*��l���@>w��-T����bp]U�[�_ހ��w�]����G��î��t���ܲ�D����߄%��C�^|�{v��S�qŜ�Rp�w��m�l��v�e����h��{����Û�+{��1��O\�j�ya�˨ϸO[ZOާ��4Nc����ܭ�^`�[܄m��0MMQ��I%�_�8�CC�)1�N�$�`��0C��E�T#퓠(�&ASt�Ēl�c�c������^�L�P+��|��������64�D r�~`�����Dȅ�߶��K*�2�s���A�,/�:G!:���TW��C���FFV6�北"q,�h���&N[f��C"q)�
_��H��.�����̀��vUO�a�������L}Д�.7�ݓ�C��D�;�Ay�L�'GYw�b�ϼ�lq�a�}�΅ ٠�Q�g!��33�"�k�G����(�o��Ӹ�չ�=��](��#kV3끶�Os���?��![��O-��<-�j�/�^�v��	� ��n4�f�����]=�n�k6f�x���M���R_bM�. ���X�{*�ۂ&i}�A�Q�rհIms�Q�H�k{v��޹�;(��5���K�[�TG[/w��v��}o�Mk�1N�Z�<� S��d?�(m�}+���GL�͌�9N�j��v�Qn�;�ᐃ��-"�����j�+�VR��V�om�&���v¢���~��Ԕ��,�w�a��Ղ�JxR�{��gdϊh��&��R��$�?�Q�����s,��-�ޝ��������)�o�'ǵ��Х��q���@r�� ��a��I�X�$b��F�~��<I�yw���`% ��$z�8?.��o$����ު���)�<F�覝��Mk�/�s�E��'��������d��ɵ�E�3���m�����&��q��͹b��Lγ���6�o��{��$���q
��
�P@S�����rB��	��,��Ī�럿l0��բS����p��Ҽ�Nѯ�_F�&�^-7�а�4�M���$�������j�czWxP-���ƶ��[��
�Ȋ�w0z�Y�����7��G&�+�:tc�L~W3�On����-����(�g
��Fm�۲R�'|%�s�zh*(	eu�Y%Ɗ.X��$�m(���A��o��� ��?\���2#,c���]X��d�ѷ�~��n¡�����Z���t���R����C�����t]l���h�˶�NPL��������ݩ}h������p騆�3MA��|5���o�8���z�4GoͶs�E�i�����

 ��K���>mEEO�TW�T�i�o�Q�$y�rA�Rw>��iy�/�e#��r>n1�`�#�.�'Gwލ.���X�_>�uO8�D{��7$����ak�����d")E��k�ೣ:�M��rP'����*���5���wL�]���oV�hpOME����n¯�up"%�p�a{�vtge�`{=����Au���@�}�b��Hw�$�c:������4�z���z��%o�����d�k��mc����5��#uko�����ˣ1���0-�����֡��^k&g���	���e����6��伫~r/��?�W���*�I1����4�	��s9%.�������B`�%x`�_��g9��V6������y۪8�`,FsPӠ���2���<��J����Zģe��ę�+H�&�e����ط!��,�UT4�?e�<%����� ]��UcD���X0:�)6��?�^7�ٚ��5x�CP�G��VeU�����s�>�>hc���3\�J�w׋�$���O!��� ����wX���Kf�U}��� ������)�������{L�N˂?R ��"�0�o��&���4�Ƿ+��Z?��$J�1V��sp���5�s
= �(j�f��rL��;5|>L>都�wPZ�\�#+�?��X�����*?p/�_G�嬄����[G�^�,���9�����^���|6yԜ['�^� �|�[{�����Pm�rb�/݆�O67�{�?�b�����3k�5s����$��A�&A���Ĝ�O��N]p�a��b��-]q��+o�Vm�M�m�D��òf�F�q��So;o �a�҄�u��.
�\����`�w)vO��/�i\~�����F��|5[����Wm�Z���￥�q_��ρ�=x�c�thG�5eR�Yÿ���@<�K����|6#(��CS�D���\ާ��
��� )��`qт�gC���E_�PSW�e�b3�-���A0��?���p��3ͺ��A�@��b���q�� ��"�Jr��Ւz��*�L�:g���T�*�	 ����4mV�����i�� ��R^���x1�=8-M�u�V,.qaaKx�_�(�ƻ�Slލ�ЇLJ!\xm�0+N3ֽ�:�W��{5�l #v���A��GDG���z�vفtÓ��)�B�n"�I��&ް�ZR���,���n@h�[Pʈ���m�}�Lޘ���C�s��O�`bJ#-t�"�_�]�[h�d��rU����q��d�v�F�)��PM�>8���bV�j������6ۼ�}��o�c֥m0��EV�����"gfS��b?�2)`���������E%$������'�K�I�V�T�H����Oޡ�xj1�?�n��""!���Z��#����c��?̄#�-G��I��P�u;��sl<���d�ϵ��M�r?
!�/�l��'�3]]��h������a7�)�����)!�e�Uǃ`!��{QIu�g��fR�9���3��f7>	D��9(�!Z�^]�~/���S1��7���^/�7ˍ��U��)ؙ�?�#����Vڮ+�'����M�_&_C��������V|6j9�&��ûZ��Q�b�;�[����|���
#�G"�v���`	x�b# IX}���47�AI&��`Z���û�H��.�(���G1/��(nc�D=thXs8hӫ4�������[���}�*p@&��;1U�/D�_�ᠷ�j��F�Pd��t
���!���i�ML42i�z�%���+K�I(�О�so'Q?CK����c��d��o�c"�����8�y���JU���+s��Ҏ֜�"�o��T�%�]˃؊!�Ĕ�<����c,�;�������8T��Ĳ�`XJ|��4��ټP��p��&�{�b`_X�mթ�}����9���w=z%�W�������-��U
Ԥ��!�\�Y�%h��F�_�}��xW{�:��~4q)�p(i��y���x�g��b�%��	G�4�b(��ņ�~�a������h�KbN{Wzc�,@���[o"��A?φ�$����Fm#)Mk�m�1�\�*]�8s���&�ߢ���L*�����	�J�"���ɣ�|�l>:��V��*9)cl���W���l	P�0V���%9a�E�9����X��("i�E[�)Km=��&hr�lAp�R������M�����5cFau�"��&�4���n�ӗ���j�H�A��.H2m\�L�������'}Yf�YL����uݻ߂z���z��:?IeoD���U.�7甜EAU�v�v��T��/Z�Q��eD��d9���c3V�V�؛3�]��L*:$i�k���<�}L�nf��f���,�3Am�xM�b[ø�p���Uj���rfj���.���"��8e�QM���	He1���8@�B�D�By��ut��,��1Y_<��"LcE��KI=�y�@����&�-<��C�8��,ݵ'�=�2�_0�Y� �M�f�+���|�_S@� �Ɉ;��I�����5UiII��j������Z�S�����E��N+*:��� �w�c���g�x�L�c��Ԏ_��Q�ϗ�Yh��HL�h �M��7�὏�D�L����� ��Z���uk�	���H2,>�T�W�����Jy53��e44CЎ���=撎#1@y������3��ZW3�ze�ukԐ �h�Ϛ�**#�� i��"�݊���K@
��N� �}[�6M� ?LP��Ҫ���|���,#=�/�ȑF)����t��n�q����W��Sխ��q-G>�9Lq�͒�٦E�I4 	�#��r��6�W���T�A�u�ͪ���yRp��Z�w}�8���І�~���%�ij���z�h�ϖ#��NQ�h��g�2eC�V��'��9
�����4rvŜ;I��K=J�a`͢J���_���<T����d)ʋ����@��/ԃ��>F.~E�D>@�c̦�,��������-�>Ѷ����f��qUȊ&���K�>��|~}����v�����g��b�^�����Ƽ�j�)���K9�����l���a�����/��CU��N~o�"^��K�{��^���'s��:��;�+�PP?��sf��?�iO
��#��]k]�`Ţ��>��c;��}�ӳ$L[P_�#�+���3c�g�F0�G����#�6zK�(�jC�ͣ �(�	��oi�?���(:�;��X8�d�3 ��J������z��zj'd��j��1�溯jLBW�N�~�*��n5S��zȓ�ԭ�����`4[����H�yv��r�Ҝ��M{��I�FB���.�4+��Wܿ�響e�η?ߺc�ޕ��/K~4�ߌ6�g$�G)S�!c�'����`΃�ѝ��D�Y��[�2�$�툐"jH���%�.�9kQ��1~��N��#�7����~���[odf�,���`W��O_X]�*�����&��y���r�x���P�)��<M���V}�����0._U���c�B�e}�������#���ҧ^Ǐ�C��T����S&�&Mz촱 q�G���7G ������&��J �#�sDD&�h��� ����?lTOY�ٞS�9��OO�o�H���h;����mO�`'��P�Ez���b�ZwG"��M��m�j~���켛��z��>�|_ݘ�������{���}��Ψ�x�����ӧ���f��cx=�,�����e{=3��H_G��8� ���6�.Ƴ�T��ID�8Ϸ���`;f������a);�%��8O�J��JԀ����;�����E�`{5B�~|����_���B��I6�0�U�ۍ�}W������`���z�r�ݳj27"Sl��m/�p����X�ˬ,��ۡ��	�-F;Ó�
���k��*�x�<�<�|�FgB\�- ��欯���C��$
�Z�1G��V��u���q�!A��5�a���ݐ��u��S���*e����l��K�ˎ��ߋ�+��M�1����t[~x,G[��Z��΄^㙅S�\M���|�� ���5U�H�v�]���PT��#�%�⁌X�3��A!�$|e# �f8����Os�7J*����P!��95��XR ���ّ�+k�&�ߗ��!��}ϕ1MU�����K��-:���9V'm�q(�i��wc㻧ά�	)Q�G��}h�Ȱf����ߒ�S��KK)�H�u19��c��£�U�$�U�h�rL4����Y~|Թm^;(������͔��:&x��bd�bK�I|�"�"�?��[�#%�z6(��`��B0��k�:�����wB�{O7Ҋֽ×�FΦc���Ҝ& $�i��MzZ��ff�>:����CG����#48|��l~r�*�tV{�H��4���$��GZ�Zbm��㿞D�ҌrX=k�?S%�ޱw�G�l�`+b�O�W#�e��d�9CM� 
~#��m��_��6����1��v�#,����c��I�\X�vH�"x!�Av{��o�V�XK��Y�x.��_	��?r�_@��#2g�(-�oh`p:�����p�Zos�^H����$KN�?��m��ƛ�Q���k�M{F�S���"*$�m9g���|����X�<�=B�����>Z�%��}a��>-��Tw�#���f�n�՟��n��V2�,]�>�H�@'�`D�p$SV,��TQ�F�k�x��A�C�:Ԯ�USF�E��i��c�"���d����+����T6ex?���^��I�	on<��<05?����Lk%P������Ԝ���<��}�A���k��F~�=��Uپ�]�^g�nK��&0�_O�X���lLbەj"�(]k�G����c�j��H4���'l��Z�56$�}޲`D"$��F���h�u�����RlT��RC���/�����}-�,������I�Mc���h�q����V�˽��G����p���f*^��xA�y2����ˇ��e	Q�h�|!!����ʃ�6�m�,���<����e����i�x;�F�)�� l���I޵uW�a�dR��5-K��{~�E�zf2�)%����f�c�l}����6]�x4��7��	�@�U��U5���ܧ�J@��F�����`�Y���OGK�0����͝_t{����
�54f1{ؿ�p���&��[ԃ���;i��aQ��������̀�������拓�4�rxȩk:E.�\:�|��!�[]���{�� ���*�a:	�G�s��@�Y�� ~����x��\�ߥ3;7�}4}MM�bl=�����.����̠g�\ɱ��ŁBo���y��!MV_h*�z�����8��������!MW"�D�d��Ao&w![�����#�Mmac��Ca�p��HN+��U��_��o��J���+t��8"dN�!�l�����o�(����@0����"�k��P�f�d�r�sd��~�F��/O0�c$���~lZ��������Z�u�����H1�v� �<�C�T�9�Z/Z�PIJI7',�aS�uͥ�V���n;����<"we=g��_!�l�uu��R��2ι\��H喕��9����"�l��I]$�BMZi�_�_0�圝�5�9�"a�"��--N�#�!�&�oeJ'��z������s݀�rr����@������7�w늲^'e�+��z#��ci눆0��A|������m�G`4a����Pl3卩[܈P�#kٙ<���m^j����#��}�1:3���<,C�J�����-�-�,p����C.>k<=�m�~n!��DM��)Cn�9����^-��
T,	�0~=f�"���L���eo�qrd<@H`�zK�!�h��d�A�,�\ؿ���s�1{�i������W���A�1d�e[���rʅ�{IH0�R���S��V�=��^9�oRfq��V�?�� �Ȅ>UkY/��k��d��
'��-��lu�CزOb���r�y�r�)�7͌�{�Ǉ/ ��{�L�k�/P�౞�3�4k��������	ifv�A"((xzmVV���� )4�(���!v9>?R�6'���/&��׋�n���A��+Eh\%�<i[�0�qzm���˨���>�Bط`�T����づ�\-�ul�ĖF�*�����'�.Q�bi����������ۯ�^��4�f&�JJB���oz6\8����ޓ�Ц�������=��}�} ����W,��M2b�������n��˜}�*-���˽�P��,��_�^9��ZǏ��Y'�����BceE�F��{K�P.y �MG!�V�V�~��󉫷Y�|\&���u� w:� ?��Z�!����t��ָ�$A�k�SO��M-F�"��'��XD���`A\�P�����n=(Zc�wI-�1k�s�Kz�`�`D3��ʥ�e� ���vb)5���1u�	kNs��
��^m�e]83{���ƥ�U{��Qҏ��Lm��P�q>W����h��� 7�<���R��Qu��$CC��*���.S�]m���s~ܔL��|�;b3�}�_�F$���&�94yf�ۦ��y�"��7j|و��A*;����u�S���;�Xҗ�������F珧�]�-�w���m'��-%}���C"�����v�6ZW���P}f<a�Yk��r|�Fõ�n�Gѻ��t%�s)���n�hk� �>KZM�Ҹ�L9�6+ױ*k-;�p���&$�Қ�˝C��"�N�S�%�ܽ:O�𲜮oiW�J��l�8�f�Ej$z���b�?A�B���x�~>x�@��r��Q�'��b�\A���Ӽ��"�����7��
��x$]�O�o�j�����i�Z����n4$b�<8[�b�d��yT��(��;�{�M��o ��Â���1���M�X�Lckr �7	�E���NXfI�/w�
�?�h���=���D�����Z�����9B[�j�P#}�FL�~�r�G�bS�3��՗VS��1�8����Z�A��w� }��ތ0'�<V5���v�`ijjML�����8��Kv*�5��+�ڬ��P��y����Q�e\y_��L��iOg7	b��0��4@l�LLNv\�0맱��z���� :{[|@��31ǽB4�}���\\/�p"'c�g�i���Ix��^9]\^���8)"E{�}\��0r�+�+��.m� c��<���yf��F,��6�E8�
tvs���.r[�.|�DH�x� uk]�t�7r�4g��p�$m�o�Ɋ�3mx��hR�%�gw_��7��/��N�/w�'76�f��D�a���~<�����pd��{��n��X�����K?oo�����>{r� I�5��$��`��W�`I�2ߟm����F��8�אd?]F�1�9Np���
��*��c:Bh`5U�6/������^���F����3���<X�����#�%:1�� �W�i�z���b��4�^�ɣڱ~i��B��5Q���ƾ�TX)Z���m��Ùb�?�v��U��3Q����1\���|�۞G
2ĥ�$���Ԩe!�����X�b𔔤����(3�:-=q�����҉�z��Q�z4���U�	[��Л�ɓ��.�'EL�Wk��3��ۻ#�G鱢�UT~�r2�MH�Kq��n�c������e���M�8\򣬻�V�yLR[����U��|%z�PH��CDaht48�M�뇐��eIJ�!��js3.�U�L�_~"L=��݌L���u�st��Anz��Ua: �L�r�~�Yly��P�.������G�7��_��~U��M��:���e��Pu'���3��*77)N��x���e��0����~�Q��j��b>�j1�b��u}���[�֏��YK�	%�C��Ɣ��?hk��a�~��޻X��}U�S#q5��FUެ����xk6ڐ���{������z}8�㷭��������&9���M�0�;y~)����;7��d��nTռe�i]3N���O��y�������BWj��X��2�4\e�a�ݣq�@��'fI��ԛ?�wE���;�,/��<<���+��u6K�i� �?\� ��%^0,�j!ߚ�:���6
繮�1��������Ի^����c71�:�Mn�Q����F�d3i�"_CAۛ}|�턁�t�{��Kx�9> َ�,(�p�Y2�i�)ŐQ��-�"W�G�rw)�!��*u**��N.OL� ������i�bP�x���(��ei��p��m�'������{&��Zg9&��.�{=9��#�����Ū���d�us+�ݷ�M���彽=�vھ}A�B�@������J%�����x��ss�O>c�.L�j;�߳x��!���
n�� �u�*+�A!KP�#��	��]Z��I��"�Ƥ{��nnkkq�!988�MM�9�s&�(S�Y��<ì�����������K=J�ׂ�=�0��H����)��ńo�@���gN"d�%�+�gD<V��
\V�8��oћT�_Rs6�Zr{}�2�\_-q�S�m��S��A�e;1`�h�ڶ�@�Il*�9�p��6# V�3F�7��w��������CL_�,�d��������Kћw�Uzm��ˬQ�0f���djH#cN�AciA���_@��^BBB�����6\���uu7:6q�'�}���R;���g��@�[�ip��a����E����+*lR��
e҂�m��<8t�n� #��Y3�>�5�'`���H²Ň��/:gmv�1�uݦ7�],O,���$~.]J�/�{��aq]���۪�������5��k�g�f����u�x��$���oG�".5A�׼4,Й�T�*А���EUe�e�eEP���hWܐ�β�`�;o�k�8)�'��*�aK�Oн/K��J�I�5����W��������a>���������SBQ�~��i���K���f2#M�{���CFV�XT�ߝ���dҩ�#�+	vvEyy����c��lFI�td4ES��L*9�����dS>����^�������d��5@{Da�-w`?\"=���U�������۫X�U���sÚ�	�4�%N���!�|Шҭ��H�9&dƒ���!!�s:�,,:��{'��6gg����K��D����	t�o]~H����+�}o��g7C�1�b����Jg��0\�!�p�f(��ވ�q[�i����	qV+۟?���^Ff����&"���O��x�t[I���ޤR���ۑ{��2|xqY��&���췿2��2�䗖F +>#�j�3=gFݪ��ӓ���d+K�e5��@��_F�s07�2��h�q�p"�����ƛy���-|Y���	Q�:��<Ï�TH$��;O�G�,|�P~7����Q��> �g1;7f�r}D<�^��Ƹ�v�R���o3��#�^�ɿɍ��Gy@ņ��jnlo�.sg�>B>��F����������s��WڍY)9�Gm���xn��������3[�׎���X]�;vH$fJ3m@�\.Q<2����p�!-��&�d��ܣ�l���Y{�jowR1������ע寐Pܑe����dt��x���K��O�Eg��Ʀ��!I�>���0kVlղ�**
*�u���+����v�7�F��Üe��/7�pi�ץ��㦞�!�����2���I�
SRt���,��$�e��%me���<yd���D!� ��ڭM��C��5F#n�e���>d]B�M�w�Rᄴ�D�
������>�ILX���k�(�q���r�r�g۲�fie�l-TR^u����T�_is�������NDY�Q@w=�ݍQQ��乀#�-�Ǖ��x���;A3����<�^����Q[d����>�[��������o�e��6I�4R]~/�/<�[:םg����^�-6��]�Lg �^d'� ���ڒW#f?��"9r:��6���*x�����������^�1�7���M'|��'��S�	9��m��������ekӕ�av�k(�ؤ����������'��]�b���9 y��j��^М����̩]|���U3��[w����B��W�m09���H='^���ҋmF�� h��S�ǧ�6������Ԍ�Q:�'�����Yy���_)II�<q�������ٵ�K����K�S��n�f��w�cZ^@��6�8J�6ES�|�i�-CX���eSkJ�Х�=�"9�Xtz��q���̿v������	�Um,����+������5x׺<�T���I��	���/9��t׺:oS�ř�rifb�o$p�2d(h�V|^B�mn��,�Ci����~��$�bV��?;���ƹ�Q�y���W;��)�E=��
e{��U�S����kK;( ���;;���̆s����2�Ŝ�����=�J��c��t�{�p�^�� ��Ws|�X���G\ΥJ���I��/_8������׵��I��841�I����6ߞyd������-S����Q���u����z%����
!u>؂��i����7=q�:�n5zA-A]�\q�a��+aξ���T�֘=�y��5����Ӝ��{_��^��LΙ��|�����l��5(e��Or�a$� s�+(Y�XZ��1uz�q�<�v]:[7�~1M��(o���K��1�gMm6se�p�I?���L|)�G����`AB�ں4nî������4	Sӳ�
����X4#Z��l��í�*�ll_Z�*���L��^#��ם�����A��"'נp�Ec��F����L�>�N����ױ9���ډ��3\��;8�����P���7W��i෡%cɑ�q&;�ߖ���3/-�E�l�q���A��BaNE��=���5����4�c�r��/[N#�y��Ϊ�z�eP�~Cf�j�9`�^�K3ff:L�2⋑'��m�l���izތ�Ae�1U���!=������0^]�YL�M�1$��[���_Z�I��j����<�K�3�[�^3j�YݺcG^6�u[�>bZcu'������UPj���Z&[���J%��}�w[U%v��2,�Fw��\^H��'v횝��@���� �\]¤�PDO�6Al�����	U��k��,*C:nׇTk����xdϵ�f��_�q��g����\�(��ޒRy����w5��-�/�D�zN�^����b��:�H%�t�@{6���>��3֤{��$7���8
�NU�?"J�KP���:����4������mĆ�
Զ���K�Z1�bI&������JMG���|��ץ�뿅����3��*ٞP��M)<]��Jd��y��oFw�u�Q�Y^EqS�Qs�������3EU��X4�_��v1�Ip�0�4r������I�DE'�o��˥�'���@{S��Q���z��؎�P��6|)����/)~�����|��r�z��ʔ콜�M,@��8Ϫ����á���U'��}U�eM����zgV{��W�������e�߆����f��3��~��'���K���vQ�8ڞ���<�VU��ڥH�3�&�6���0i��W���j+�1��\Z��>;sh%S:B
Hq\-�TW�t�+-ݚ�{I�V��tG�Ur��+t#3|9��C)������~_SB�}{�T�>2Q 9.UԗG�� Q�r�2�K��?��4r]V��;�Lu�TN�y{Q26v_7?�����\!��WF�t=(�>W`*x��k�ۆ{#�X�j^zYt����v¤2�3?����j9�'/�5���N�{���t_���}Fe���Piv��n��Ƕ��F��#��׺��ho�����*���,P�������W�3;�!����M�v��)�����j�́@��z��>�
�Wx�,�s�1Ĩ(�«i������9PZj:����4�s����@ySH*޼�17�=���bs8�������^��K&E�5`�7;1Ѡ'�@��|_��Q=d{_�<�_̣gXR>���q�=p��C͐�W:04;��� ��u���~��?Fe�3��9�b?���������|i�9B�Q�m�I;�bg����fŚ6Ջ(���՚�:��Z�uQ��ecW��w3���Z(j��އ��l(���R��^:Gp�ȹ��4���"���m�f���z^��B� ��9��*�5�b��>*�Û̢Q��NLR3298�?�z�TV�� �:��I���
F�3t���Q���a� z��\���yƺga��~��x@�vd���@��
����Y�3����lY���J�p����@��C	��B�Nm����Ȓ�P��b�|J�Nc�4E����1�����6gx�A�Y�n��iC�{(���&�pK�Krx�u�v�B��X����"�����''ٽ�06���Rm����8%&�Mi�j��YWg�ժ����>�	����b��!��s�ޅ{N���B�������7ص�]������[F,�G�Ђ)ʰ�o�}�E��<�3`�<(����Ŷm6�cb&#���oێ�y�qqT�f��}�HN}�J���D��.�����Jo���+��#���@|R�i�r,����xp��MX4=�!������r����f����xϰ�@0z8^�_{V�~���
+�����N�i*���9�����ʺ�b���I��0'���t�	"`�r���U�ol�Y��mop#�J�K��G"���k��� �u,�d�����������vmu^}�r���� Dzl�@�� -��L�+G�Lk홅��x�)�.�Ԋp]Q���	�J�������i���s̕i0�T���"��*�M��d.�uE�,��,cj����B���rP0��k0��Ѵt%����^��?	?���I٧B�����#ń�
���оt~�;�����bz���oRS�ؗ��sU��q�����i��bP̴=�f��1Uذ�B@�#����)��b�K�(|cSmQc�����4��H�?	AI$�	�v�����M���ľ��M��<}Yz}N�1�ƻ1a|�:�ٹ�Zz��PҀ��)����S���l;C}���x�>�r�p5��Vba�Q� '�qB�җaZ��Y���ʲ���Af΀�7�7*��@op�7�9Z(�wa�)ǕV��*b+�-M���#�^5KQ�A�Kz���x��?����|�p�
��ܳk03*�"qm�^k�^���sہHqT&��Jh�@��ߨ�����y�[e��4_�$��J@������'�iH<"����ti�ѿ�}�ӅĨ�z^0Z�'%G�"R�/���c,>
������̲�fx�\�����n�_�Ș�f���`��^�ϪT�{eO�R F��C�/�����o�Ґs?{��,��I��:�=�����_��
�6�w�O ^�f��>�y�W����شCJ)P��������-j��jNKJe+��,,f�4����-}��g`�Iy�,�Eg=7&q癹7�W���[Pd;�Z���I����⬜�mjU�Sa��j�h�س�/�7lاN��6�M{5�6�J(�#��/y_b	;b�*���\�y�����J�]?,���_D��w
���$�i?i�E�������D뇗�'ZN6/��꙳����.��g��V٤�,J�3E/�"=�~�3�i���O�<�z�_���J'JM�G����E���rb�>��4�M�ip�uu���r^�q+���i11��#xU1'�Y�	�~��h�z<�m
�o�r���1B$I��i~u�$�����&oy.K��������j벬���.����D��憒�h��T(���n��'�Db�9R.>~<}����JB4i��<��׭�|�aR���.����--���Z/��c�G�н�xs�W��֑.�����4����0�A�|<c��c�-��?:�8y�s^�xyF��r]���6@��{}Zg�ǳS���c���������F����fC��XB������[eg���#侹�dJ�TMR��lz�!;�ǖ��Q��2��P��ʚ�q0�p���ӝ���q�t��U�	Qx�}�^���#��K/5[B�����_�w��?:��Gޖ�}e8����3=�� 9���Y��-Og�˘��*J(�lD�
^�@���y5ɣ��R�����a�Z�&�׬[&���s���A�sՋ�&��m�
ԙp��46c����^(�ٗ��I�rS!#� �??����,�������-n&wNr��v]����>;����SW�mi�{����?���Z���ĳҡ�NVB/z\�*��;���� ���r���q��N�{<��k�|gQ!�c��E��h5]�J�<�n7˙SGk̷�"��z|%�5�0��v���8R��T����R�G�z�?%d�I��aG
�q\D'B���߆?���`<���0�0�쥅6f.h5��,uΥe�b���C�{�S+�\�Ԉe�,����.����$�Wj���VJ-b�!�R����F��9�2��ӎ3���p <?�z.mTP�U���PHnVA�� �?$Fi��°�����yR�J.:3�`3i-�GP9�����?�9:��{�Qc5Ic76&v�X�m7��ضm۶��j8��w�|��Z3���s�u}�=���{���Aw��!r8�}$\L���ԛ�����A��������ޛ?���HU�&����0��$B�� =�=�
>g2-r��5�0�??b��T�^R�y�x�2z	���}���k��1:�	�)��-��`5�R.���!_�$qBud�X�
b�L��xL����2,C��4�'6�_'h�/�����Q�><̡� fd����h�� ��~>do?(�;2p�L�	���x\D'���h\k�5esZok7)+�(:�˛!GυB5�l�灝�*�S�[�KC�����j�!�ڣ�����{��z���E��}��h���n?�7�y}��=N���t�(-�������w+���#|?�R:tY=I|�V]֔���ܲ%� F�Fϟ���Q�#! �K>�=Lw�&��3�1z=����p�ބ!�������g�bH���O�q�<���7>���x	�y�TC�� '�v Y>��]�wR�s�Q�s��h��n�~���{�h��ˉ�����x�H�뮑��t��Mm��W�q T��N��C�)+-��A�x��64?�%���_��Uh�ݬ8�����fPb�(�b�����k Ѧ��H������{�j�^��gaj��I��у�DA�{��%/�V#Ԝ}<u�o�3YؚV���w��L`f�P�B1�DS�#K�k%'��d���|�=�O���X����3���������qIS�� Gy�@I���so��n���򸟍��`�8��)��.���l/V	����u=<6��*�ɀպ#�����k�i1[Z���|�$pAb��2j�F�k��h�}` ��[���i[�sA�pqd��t{��[�.Ů|A�g�L8Vmá��̒�H�{*����'��8���ݣ�T�P��d}Sì�.�Y�HG��چۥ^O2�i�m)��_���-$$�,�������N����SԈ�_5��KdN�}�PBI��.Ѳk�U�����W׷#��ϧ���4-@#��XNu;��{Hթ�C'�c׽�v��B�b�,�W����IP�I�E��q�Vk�s��OD���[���L̡\�2�M�.F>3�0d�@�L}uԵ}�OJTA7�Es%�V�d0��5��A�y� �l���Q>usf��e�>�\i��$�JTDA���,#-<6@����@�SFɓ֦���bI"V<��^��E���l�-*�W��H�&&�Q�&�#,x�Tvʩ�Ռ���4+�P͋���dc9J��΢
9��b!ׯ���Z��s�h�Zf҅3��a3��i�ɩ&c�d��Գ���JQkJ�H[*�X��^_���F��H0�8a~"AOg�4u4��[l\;���8W��S��J�:"�>�&��l���E��]7LL�v`{�1��%����0֙K��H	io�z��<q�g����x[Z��dr�-�b�prwqU���ZVB�k��YY�a���$iq�ʡ�AMTǳ��ڹ0�U?�gh�����
A�ܼ,*��+��)�no��r��I9���Z	wt3���2��_�D�?dj����!]���S�ߡ�(��3lF��B����]���η�m��H}7�hI�Z�|p �z�p�tOfQ��n�y�����K�@'Fr:yO����ٌfl�e���f�[���K#K��aϥ����4��5�F����$RaD��`Ci������?_77��]�#����et�D;-�h��<p���l�XD)�xFa}#���*7����?��!j��(���B|G�$�ʋ|Yx@���Bs�9	fx'�l)r��Q�_מD7U�iL����`X�]56*vt��iy�L���jT��9�����{�|�	�>X�� -��P�Un�Zpt��F'��^?VK[��Ǧ.]}7o뻺����a8�����9�*�r��D���x���램���n���m�Y��Ө�>��=��W��,���!�itf���˘��Wg�L)w���SzC����=N�V�6�FJ�Q��R˦Ş���Y*�O�,�v�X(g�7�Oe��o/	9��r�N�:KA�(�0_����aOv%�cc<��2�����R�Y�,X�9�I��p�e����9�{
�*�� +Z|�d9�iG"�#m=ro�(��Dp�Oe��/��")�8:
t���$�/Cy^9�4�hI��IǷq��1"���r5��� Ʀ$����y�؟CjleK8k!|>�y�x���a�a�����_|}yO֋�䨢��LU�4��(\y��8��t��u6kRv��>����f����b�|QV���b��Z����.�DIK�x�ֵ��6��ܜ�#�sc�9�ՐK4�H�д�����i���4ɤ��單u-\8����u"���ԈO�G�W\]�E�m��W�_r��=�z���f	�-�˃�ѕ�a�ߕ�7(����?^����(�q3�l��l�k:Z��8���;�+#�W)�[��zj
�)�<�����u�{k�����?c+ߚȢ����y�(�89�c:��1~Z���d�d� �:�*bG��w����* .b�s@��*c�R��d��;�38�\��"�@�[vO�&�G������O/���W_a�![	V���4�Cq��GҶS��+t
 ��̐��׎��9��S�C�����#I��ٞP�W� ZE�g�	�'G=i�̈:�g�χ	�==����-�nq&�Á򾱈��K�*(?!}@P{����4�����g�]�~P-66�k���������#R���Z��@���o���0�����}$��˽���u�y�}n�� 1"	�$�K�t]p9�tں��P_q�Cu�;��@t�2#� G(�y��6b|��)9�f���^NZ�(�5��E������]�1a���|0tę3������00�3Y��JR�]�vz���λ/�P�&�P!�A�'XolpL��C �"�5�\��ݹ������F"�.��� Z�9����pS�+L��N�4��#ui-�k#��l���O��������$N10Uy�C�W��7������S鉦��'$.�?Wg)�|ō�Er�=�� �C��g~���C�.��������n�p1�i\)���=Q���u��0���~B
�Z���G��Kwg�>2FZ�jow�3�*�ɨ�����&���CG����'��'^Ec3����y?7��9#�'��G/�
^=��?yKVd��l�뜔j���vP�>S���m��n�W���[?Y�vP6�`IA�u���s[��/����T�`ꭓ��#_�B�z�6[��CGCN��{?[vٽ���L&��̓'`���
����^VGf�>E#��4!"�z�C��̙Pp�U27s�N�P�����Ǫ�Έ���Hu/ �;U`���y�Uu*s���$�y�zk���Wk�2 ����M<���#p+6�9=��_)}l3b������*_�� ��a��D�0T
�i��r�.O�<�nh�3q�f�s1�-3F^��Q�����[�s]�Uz���O���wV������.��F��U<]کC1�Ղ葁m'}��W�!�Z.��9���.��Me�u$���5H5����|ʇq���N� *t�{u�/T�����n:�b�h_��`ZR�T���5�XK>��U�f�K�U��1�~���7�Ҵ{�5[+��u��ę#A[�'A�/δ�%$�DaMb.�2�~G�|J�yi}�ɿ����F0ic.�C��O��^��W�e;���3d:���R��`�|6��8��E�*��%ɻM$;a�����e��w �����ng��&�>c��>�0v��@�X0(�H2xdƑ��8��r�=�=���IT<�o^�}�)apa�&^��������cd: &c���n�}��-S���uL�\�u��P��E��'���MTL���h/҄2?��m}��ܼ���g��0�X��IچdjE+m�9"��120�"��Y���F���[����%�wR�#ș�$�2p�.Ǆ6���Y��h��VV]|>��{�1��:����i�i�������>��a&����s�G��=��i�t��֞7L'TA��ힼ�����9Ҫ�9���*�?1�pD+'L�;�����ֳ��i^�`s��J**�T�F,�x3W.���^O\L<Ղ:K���b�G�)�ַ���n�s�ʊ�vCZ�lI�^���@V���U֫��9U%yq��;T���q��N��)F1��*$x2�i�/��:�\ܑ%
��)'X�`C�?] �\��ؔ��]�DJ�lY�]ҭlݙG�-\n��<�?$#|%J��������=Q���s��|�㵷wڂ@����T�ݫr�s���r��K��ǡ�p�|�"���#��1j-l�^�+�@(��q�H'Ośh�H��y����g�T��fZ�����iJ��m�����~B�"��i��'�+0&��Nl ��?bf�R�K�lfvp��� ,N��bܞ�D���KM��S%�U�P¨K��s
 ���{;S��N�I��<&�~.��[�,>�f�Fnn�Y��e������奯z�ل���%Ŏ#��3d�㺞��p���C�c�6%��\���/��4N�"RQ����V��@)������v��;C*4!qq.S٠Atk� s��?N:�u����W+B���9>2��s�vK,�m��M�=�a_�Ek���H޷�������p�P��u�@li�d��[%$-�#h��/�ГZUc�~2�a���P����@���aN�t��5���}�{o�l�a�ބ�N�F_]v�%¿��q�WV:�{7n��{,�]�B�`ӼJ������t�ώ����u����	k�9�d��6I-���azB�����!�P��Q��������9������#<��7���^��Ǻ���JʲA�2����z��h��nH�KH6`ʰ�~o*j���A%��ujs$����'v{��j:	�?��p:.3��]õ�j�p�^�##�O܋֬e��m﷽�ʴ�Њ��͇+ۑE,���|0Z��J�^*[�@lTQ�T}�+�	9i���Coe��G�hq�_(�ԕ(�<�=�3��0*'�!���Wb��i�/L�fy��V��`{P=�u*}��D7J=H __S�Z�q���>k�K��7<�X�^�S)�������Rr�K]c�|���m����3�GG��V�J���^���s?�p�XM�u���/-uV[P���ө�j����d��sokz�t\�MNzU'��=�7y�eY�L�ݗߑ�5)�t�a���S]���nP�)߰�t��S���x6�������X���;�A���p�ټ�����ڤ��*�ʅ�Z�G��Q����PzZc�F�q�C¥7�4��z��`�Fu�Uh����.̵h����4�|��Tˈ���Sa)�I���\�;SK�W!�����NO�^�m⣳;9<x�!�I��2��
���ͧБ�/����'�:�}3ذ�^=wq�{�)�������t(ӌIk��LV-VWc�+�@�F�u�I�����_�� {9���8�(�}�7a��h��$h�
z�!a�L&go�4�j����,e�a_�A5Wk�w�e��ɠ�rag��+�|�$	:��K(��рz�f�H�j�J@D\�Fg�%�=�ȈH�܅[V+o�t����Px��><|�Y��-��M��Qr�������IC��!�ODZ����	��
�h�_�|����[�#�Q�}��yxH�g�=)������}�{Y���e|�� ����7H�C�`��a�x�Z�D �ٛs~ U8�%��;]��6p��]���S���R:��c�8�π���G�䢙Q�:��s�qVS|�Y6����1��v���|Z~N�`6w���#bx��FQW� �[V8Q���a_�u}=�N�I�<�,p"),��ч��$ �������$��Dq�e���/��*��Š^��R6ھ���m�R�DI�)��n+�T�\u�/y\ ��T�StL����[E�Я=x�h���`;wo���U�`'%t�������>�,h_�_�4�w�M^�=��ϲ�a�1`ւp:���L�_����)L�*�MH�]�E����v�O��K�UX]����^,�H�����ٴ ���!�sv0?�Ͱ
�j8E��6��+hxL�h��{���j��t�J��KY.��<  �*-��r��Grr�ل��9)K�s1��Lں�U]��}i��t.׃�O&Z��A �!u�.B�̃=An���#��R\��(N���9 ��fx���p�Vt&~&W�4#3��� z��Ip[�8�3˵�I6
d��r�1��2�p�z�Ͼ�-�Ɨ���ĺ��L�L՛�91�K��5�����R���GR�f,�*�)T���l�����B�qw�� RT��a����֬=�Ö�F�
��E ��!�G�F�c��=s�:��}��OC�t��>����պ4��;�6����`�ƊE$���@Pc	��ƐBĺ��e����an5�#]���H^�h���it�\Ir133u5s5�8s~�d5��Pʾ�޾ԫ.9=�������jZ�d��������B�c�%��b_'3J�z���ذ�3�ˇ~x8
��J`i�$�P����g�Պ�!�-$�-9<&���/Zx�֎��`��7����`�7��S1GWJ3d��3�z���<\ɛ8���9��`�r�n3;8�\��]v��*�|S0��TLI�2T	Q��iWGG��d�� �<tI�QU�9�$�.�"���'ោ�g��`���+�u8�(!G�?�G�m�~�6�|aT��+>�+~��ƈc��î5��TǪ���I�!�+55��u��1'����#���a�&�^Ԉ�� �����>��5��힨�������3m����?h��S��^::����#D%�L��-l��^���氁v�)��,)���c]��d��$8���M�L˛��p\mk�x���\Y�9���#�O���� NF�k^�lʮ=w�[�O�-/˭W�d]Q"W������9�W��q}[��V�v��Q��lo�/A����HWOeߵ[�d�t����Җg��o��v�<�3Z;g�[�W:�����]7�U
HP�IPI��,�]�T ��U�����c`:�wr��K_N��x� ��2�^v,��_�*�:i��)�6w�[�l��[@��W(���X��p��ϣ��8��@�g���Te8`�ky�Q�ѩp�%v���Y<h�v ~�Z'o:Y����rܗV���C��"��]W�z%l'��W�e�cE�'M��T��u?Y\x��^w�����'$H�E�1�c>Oӷ'Ta�W>&�`�i�PSE��9!U��T�VFR�t�g�x̮� m==��<�)�8���37�?e�8w��DoW��-!��p�(�/�Y�m��oy;x�XGܮ����m�3LA�8�@���k^�Ob,���&�� �t"Z���p%�����;t�u��ζ���xZ:�$���]�0�Ds�0��F�rjx�ﲕ��y�yl��V��P�U�>�5�-g�{C�����<8ϤFz��O��y鰉�������"3�չ}!�JPҬQ�/���TU��ccI�d�uъ�C��Ȱ�q�͙A	���ErCYETm�1�@Fg�O	�������:��	�����X�(^�F��ރ�A�d���a;m��b���s�gu%��AN���غm��ܬ^���n89�[3ʻA�ZVA���e=��s��1
)�� �ĭ��5��y?���k>��mNdu�S������3�4,�a�:���2��q&@橯�;T��z?y��E0�z��T���[�1��';�\ָ�sAڊ;[z�P��T��D����p׃���BCF�R?JVo�X��g��a�,Y}�P�@^�̼�U"��_����=/�ZgՈM��?n�I�Vbv;���W��7�M����L��_0s)�u�ϥ����NQNX��Լ"����C!���ˠ��yT/����F�`�G鬗���;�(��*?����.�n����d!$]��&\��V���I���o���bH��D�
�6�$EΨh^=��d��!{/wp�Zk�(�'�ߋ���7�ڞ�������np�r�R-e4����:��BbyR����nf>���u��%��jS�UO��V^��X��Q�lld����f�j��r�ڬ��#�c�$#[��!o�/\�}�"�����ŨS���e����Q���͚�$���O�>}���.����Y2^�@�b��<y��Nkl���0�~_8�c�(
j�*
��L!�(4�Ӥ�nC �R�'��
�ؗ�����~���p���߽2��m���� �q%��$,4����ֱs�w��n����Y�L�੗�6���P���:���1��fR�����L��b���5�*k�Vt���@�Z��� �CN���|�l������YnI;dT�̼��J��=8�P3V�z�~~�>�_a~D�np��V{��������~�Fo,�J��-��|��'i�n�-����icJ>�k(Cc�%�_Me�OT�u�H�q��n�e�x�_޻�LZ�/�f�nn1��ut3P��P��e�K���(s�龞_���)�B��c��q�@!] u��=3�	;c������'{�\s�w�=\m���cq}�Q��W�?��E�J�1�|�m̂cZ�D�J怣�=�Z[Ä(Q�tnYm`m	S�)�;u���E&9N	����$�DFcG��4��ʛe�Dl�l[�2 L�4��pP.e,��}��8�7�v����<�s�eC=�q�0B�����c�����ּ-���\��sȴɉ�9��	g��	�%�<�~6���qN*"�,����Z��Y^��p[æ&��Tp�W|\V��	�Q[�C��գ�ԛRw�:(y������w���i�)����N��osz�{>��|J>��d�.k�C�H�1O�7��V��@��7�ji���α�/��V�%DN}ב���Xl����=Ix|�P�.g4��)���0�L���6m�:�}׾7)^�s�٪Dą��#g���3${���.��ǳ��ſ�q��c&�m:lt�\vd�p�ih�[�۶�J_DT��M�fZ�9�#a����V�X��Ne�h�+�aHs�ߍ��Q����5\կ�z�=j6ױ�e���d��L��؎%))���6�[k�M���{R \6ev����	m��T5jH�.i_4＆#u#�ɐ&�e��ޤiG�R4Ѱ��<u���,�F�&����Þ �d}���hgp�Z\h�2�8͆�$G��c��o��ۣ5[_�}������U�e�-���Ɏ��T��gs_�9ޞ�����y��]�i�(�����F�ZE�58e����Iƪ�t�$�g,q1���*����k�jS1jэ�hu��_.�es�s0+�y�Lk4��
k�+VP�rtnA�$E���ˌ����ЏN�5��B@�<d��B7NZ��}!56ّY'��l�\0��ѻ8G�`I�DBP��-8c�k��N���4����PRzg�7��тK�5���#�`�-�M	�ZŴ1b��\�׼ڼ�i9�8YӼ�?�C`���}�x�7��?KA��LA���H{jR��lZ���-��Rr0�A�~��n���Y틤z*��dJ^���L���������ļc􀱅6���N,��E��	.�'�0]��17�3R!}�9׎��ps�k]�u��m���=��y�U��Þ�@����d�h���d<�$k-��ɒd���äʛE>ΔBM��4m�^���٩�o�ő�����K4*�>'����g��yeĜ3��]c�%F"?X�⊎��Hk�C�)��W��¨,h}��f��?��֊z���m�׀af�;�]��}=G.�b��FAL&Y��o� a�%���QJ&y���O�VS]Ոt�\h�V��|�G*7���PIoГs�SG�3�@rr	=&��A���b��Xv�� Ȓ�w߹�EbL�!�R{�D�u7ň���	��͑�1�J'���d}O��s�T��5����c\�A"�����8�Po����"h���?����DN�A�m�cq9�F,/W��T��/Q~-�$�J"��2sb�͎-�q9�G��Q�r &���}��*��=|�~�>t�8_f�j�+J��� ���y�
�����{e�F�~"�=�fH�6|��z�'��r[5�~�-%���uF�D�N�.7��N�^;(NBc�Qn��Tw��������.ٹd��g����Sc;z0��ݿJ<��ۇg3��.�����&��)3��������-�e�38+Y�����]>�e�jݨ՛e����S��4yv~Ɔ���fNσ�2�8h����-��Sjs����)�� ��� W�9,~�k �d� �8 �^����y۟q	!O�a@�@AE4[���F�᷉��&4�ǃ�(V#���̹G������'RK�t�I~�k�,�(0���5��m76I�xȀ�	��ɛ%R���W@[��.��g9�N�j��C�8d�׷ߌ	m$�����5��C�:̣t�ѻ8!�$�8)�t�.4QlD���P�erts[�*�j��:��xj)�}c�n�ŷ\9�w�S��u�d�������>T�U�CS�=?�e�V�dp��~��/�*�()bh�$�Y�M����}�,��.�#"��{R��v��|��r0p��ҩ�FXg��~��Q�Y�o=7�Γ�f߼��*�.j� �87��j��g�ׁK�`p�o,�E�Nˇ�'�nS뵾�{�ש�ʦB��v�]�=�`�̢��>��߿ڮ���tq�/ �rn���"Eє`��|�?�¥{�Fm��4�E&&�������!�R"n�O��:.;2��o���}���o��v_E�Hh"Xj���d Β��k�Ǖ7vT���*��C�O�Wv���gw��4�����VR��i�BA�v��T����F�I�2V�}�W�&��-pM=@�&H�1��f���AC4�h�0$Q�1������bH��^w���T�t*���`�j�%��m$��&��q؎ �tƢ1�\u�5�>�o�rț6�>���Z��-�t�N8��}�Xh��8L�"��h�$ΉND��1���};Y�u��q@������2��M!�$�O�Lj�r*�:�.�,fѺ�)�x��/��뺲�r$�w���|[>��@gz�ק����W��@m���~�FA���ޞ��#���v�,v$�NØy��Խ ���d�,��ic{+������H��C�T���8偓ݘ�����r��fC��왾��&6=���B��jƞ�yj�YNEw���2qo��O(�Eo�r�/�h/y�+/���c҆�>�i�\�^�M�d.u�G��'�4��{Ԟi���xN�|���M)l��0�
��i�&���پ��X���lgrc��#B3E\PO��2T�&�t���E0�~�/��L������Y��\���~I�O�ܟ�<�s�A��zc�Ri�op�a��-�$7�S��]v�PoJ���0��� l�!����:������k��N;���Ot�WL>��^��$	��L��4����}����I�8$�X�E����2��v�3w3(]�2O��m���G ޵�u���o	���|,�)�v���3�[�oʹL�YJuB�i�]:`)Zf�L�<�m�֗0f
>�l{+b�qq�'��h��>; d���`t��H�u�{����{�Oc]��C���a�V�s��81��`)3c�/� ������-�d�����+��\s������Y�F��`a�`���d�����n���o69L|&iص^����� `�4��5�d�E�� ����'4�͢	�8����}�Z�:�/�>]�7�WfL��2���+�M�k����HlZM�8���N�����.�H�ǵ]sM�t2j3��:�S�yq�e�ʩ Pb��)JŚB�i��TPd	�ڮ1�)�_-zKN����\}R>^b���I�&`|��.q��2�td�/�I+V)P
���$3YI�D�TB��]�\�Ǥ$��� �}�6��gH~���|x�2c\W��>A�����N�W$���#B�ږ�O0����1��M��6'�T�Zͨ���R<�7�Vo"�!�YD`q�*���Lg�YW�L������':qG)�/睷�Xm�F,w%�ָQ��|� ��ج�&}��b�![�hԉ7+;�h>Vƈ��uuWBh/�w�E��L�$*�ȋA>;���v-�ѕC��HbR�iA����m�?)U�&rh��r�)����032���}���%T?1�u�F�M5�͜|?�n��`f>�^��(솥�"�_�Yg:Ÿ�S�_��
������>RzrzNN8L����ܺ�b�q栙�J(@�ݷ��4�FVF5�\��� �ޘ��6803��8�$��\�~_<6e�*����j�Ml�cL�9$�����j:.G�fM����3������m�Q��|�OZ��e��\�Bu��_~��vzʖϵ��r��20;��Zyc�$�6jz�SV�L(#�PDi�EG�r��������s�yʏ�'�Hԯ�,�"݋�Ν�ϰY��W�W��YM{z>b��1����q�ï4�"�́��3��(V�c0;Dgh��`@�][6�X��h�*�G����@�>��g���n���n����������"�o-��CɒD�At�"6)_��uy��?�#�o�Kt�/le�꺰n�a��FnO�]w#D²2Z���z�����Z���F*��-)�-�?g��!��������Zg��fy��E��%�������U��M5m�p�ޞ�~eevhZ%�nLXb��@b�O��C�3�+,7���tfR���&������'V�fi����X�j�if90P�}W�WA"P'��}ĦL~����s����p�v��c��`��-�EZ�tZ��
U��>������.	N�k
��5���I#������=%����,�K�f�30�,�ђ�&��T�̂���P�`C�1�ϸ���L��h�ke� ˖�O�Yq�e�Oɏ��B�K����,�^Hw�Β^��M��`E��D���:��z��h�#�U`x���Ơ�w����ɖ��J�}�9#{�����,h	@�G��V��L|��,C�[�����yV9����ol�m�5eh�@��p�J^nyTVnY�]5�J�����34k�'Y��nA �/N���;�!����$�b���io2�X-���sZ�9%K>a�v��g�J}�҃0��+m{�Et�z�z���b.�����T�r����=c�\qC�}R�t��vޑ�m=�w�`�.���q#3"9�:=2{��'�8o�-�M����(�.>z�L2�A�0X멺�F�z���������l���������Dift�UX0G�->�T�z4$���`'}��|޿�D������G�iJ�,�����
Ш�1��-��f�XJCS�yC�x���3�:���.���h��8�(vSkSooIX�Ӟw�~>C�ά' q�ɕ���*���P��b�Z�p7\ ڃ��tH`� cqÕ �H+���r�F0s�!��=�_�,7:Z���h���u��dAR�-Sj�H��q��h�|�{����_��:Ri�L�V�'�@R���/�����|
)��/��0:�m@�˹��q˖�/p��]�ҹ=V1��og<rk�8��p{$�pq��`�u%u���^r�������m|5�PS���zE�[�����k�g��Q�Ze�Y���t�*~H�,��[�Z��OB�	
Kl7t�g7᫅���eH���(QȻ�|*��"G��|害L�)���E����M��w`��ܪ������\b K��f��Fl񚗐��ǣ����H?Ş�_ے���(�%Q&v��>^�ڣ���Wv��J�Zb��=�R��̪�f�uy|K����.�xy�_q��Ri�8o �ԟ_l�Q*qb���O�'�' �^����MJ�v;ה����_��2��$+��W��9W�u�/K�7u�67�MR`|����JMǖo��,�V$���$:��5C3�� b.����|����T�,m�Ym�-�N՞V��5�e���!ҁyI��T�$:#8�G�.f˷�³�'GR>�g�k�dNA�8XT�������Պ�Ez73����~�C-����a�P'�.�`xZ��+j.��e���,�����c��zl�K���Y�*H���죂�/����1���[�?�#��v���Ͱ͉>�ANg>��Q|�M�9BD*���댢�}\�樂�YVHo�����6�U�]�z����w{��r ��l'"��*z�̝�S�c��MS�o��h:p�u��I3�c�⛨+š��̲��i|�։N��ֳ�NV�#Eϻ�a~-k���O�m�����4�-�^�'��C��2J��Ŋ�D8�����cm3�o���e�l����9'��a/��p��%��o�Qh������K���f���r�~����K�������aWq]ȕr[j��
�Huۤ���$�	����t���[�-�bO9J���W�P����_WX?��Q��p5��F���B��ˎ_7�i{+���u�Wy��4�:��⺫�EOO�����KCO2VG����7�M����S��Vv��XS���I%�!-E�ޖ�yA/	�M�,�o?���4w�p�ۃ��G�Dxk<��� A�o��*� y�OP����pp¸5�R\�(��gn��;��°h.���/y��e�P�Dzo.c�D��1%��]Ȓ�ӌ�/��Kmͺc;�*a�y�Ifb�=��{f����C�$(�u����-�z��/O7j`�z��(�-�����7I�_��� (�d�0 �U�l��&�FϜ��!o*T�	�q{�<m��9�������mG߇�+�뫮�KR�n��~yla�9l���JL�T�V�K2�!k_�ASXXj{4�����t�U-̀s���u��;J��;��s�n�FD�:MJ�tD�#
\
�ixV��p-��$�&Y��fSމ6�g8�2�2�Jlw�d��ΥnED�L����J��~�9 ���I�2A�V2\�G�JDzg�n�D�&��G�(s��^�L9��f�#5LVU|+�L(�0��g��,�[��d8͗���,��]t?[��_��G�<q�g����So3�l�%��������OӬ1��M�*��Օ���_��>�/�T*�1Hο��J)f�/%�h�ih"���E6�$U����$UQ�/�DC�<.���k3=��B��O�8��;�5�Z�'g����)�1�1!C�.7�"m���}+yU�㹤Lu�;{kF�}��9��%�E2�����}��O�:�4��}o=e�@�<���K��,��Wq�:�k��h��_��_��u���I�L66=�8���.l|0�*���'�*ES������
A �p#L?H�����;k�D4�O}l5����mz�|�:�O���W�/2Ȟ�P��ߍ�=%�}���M��p�+���Ƹ�P�}�<�h�y	/�s:-��,��65C��47#�2�4C��J4q��Cr�ޚ�V�㤒�)���!�I*����D�e
���1�y����<N� ����8��p2{��`��g\-�'��� ����O##�Ҝ����m�|������Ef� ���������Qx�.Ǹ����j1
�^�oMߞ�$�TXyھ�4^�'N؁�`g�1���-Z��%f�t����*��^�I����_h���Ј��6�{�y��|U��qGp�&��#��!����7�N�X��RVc�Η½���E�`��0j�Y��74�ƞ�;h$�$���p�����۹�?ݟ��k��)�=2%7]�u��|�v�-g,�G���ڒ�����F-�j�_B��~ դ�<?T����k ���k*c��TH�YŐvs���L)ޒe��=~���[Δe0��=���է�q���\��CP�H�'xIeB��Є%�ăeJLTH�ט�	%��+Y�0m����[o��SB��V���@}�v��N����6��T�<m�p�����k��G��=�mo9���zc�ўy�� ş�����7��Uj	��Tk�q��w\y��E=�q3I�>��Vi�uJxk��jVI
zqV��L~��wg��V�,:���Y&��ꩃ��׈���
�
&~ݣi��jf,��c�������}�iI$�����D�A:��ABJ��Fb��nV���ݥ{�~��~~����>3s�癹�g�y�9��{h{b�y��R��M0m����q�b�\R�+�mC�h�ܞ�j��~���[�h�ȴ��*���qB�����X/!�)s0����-�5��y�b")�P���lp����8�8��Qt�U_
Z5a%s�Ɖ�����:<F�ݖ1��w���]���[�+2��sΏ�w�'dJ�
 �w4���B/Zo­ߙ�xt�LS�`���=)t��S7GD��Z�6	qgӶ6+�t2D��X�9�c?���l��H+�룮[')M ����ɏ��^Q��<͆�X�|�dk ["|%f�hjaZ�I���<����j�T�)�~�-D�I�kƬ�ܥ�޼Ƹ}x\�C�| �/���<��0>1�XV�6��q��J��kԍ)\��wh�;�Vh�Z@�D�KZs" *�c��.Y�+�ÿ����W��R������1�E��=��ޟ����P��!������y1�9G�Sh��uqRFU��C����uq�������rhY z���_��� �9c������]vf�`���v�}���xE&~z'�@L���AIȒ���qn���/�*��E�����f:`�B؛Dg�V�B��2<UFu���|����ODRQ�ŗ�n�f-	���!����;�Mj��x���h�����E3p�Z� ��{�-��X�O�qw��a؛(T�xA��c�I5��5��W/����u8��;��ޱW�"��j�����09p�vum0�G�ΣpZ2��;��31{h�W)��C�r�z\�^ȥ�.��~����w��X��z	����-1����L6��0���F+1[�@����Z����G�7��B��%Ƒ��A�j����@<��!"5D�jm���C��c�h�e^�m�'oa��;9���nˋ,�-'dEp~"i㉓�*��l^�I�M�]�z)��ij�A����X�j�~���c��>hM>�����Y�����<��?p6�8�Ui� ����9�D�J�'l���Ԑ->��1�5豸,��#jm�����,��~Qn,%�]	��2^���¹���� T�\{I��nQa���Ë3���OO<�-��oވ��E&N��YuF#�3����,�[�~��so>���2N����G,蒮L<h=цt�nh�~oYl�Y'ܥF��/x�����"6�|V.����a�R筁��µ���l� X�Noz�g�'Z�{����ba�.�.��Z�󟑒Wx$6>�rs���E�^�}2t)Wې_�k��3=�I���WM�w~���|e$N�z�x�
؎ކtg�؊�'�r<Z�� [��_��5��}�jcw~��~h�җ���M���~�"/��QwO�[2��v��̥��s��l��R����)��׹Ƹ�Ql���b��q�iR�`f��h��6d��L�\����:҂AILc!�0D����Y�����T\Y���T��>� E7z�^��Y�4I�)m#�l�=���t�� �	Α��K�X��N��}�n%�l��ER��g����W�j��,����S}���'��Y�B2�#E}賈�R�9�?�(�}���Ȍ2x�,Ë�A��x�Մ��ʖ��nAʑmC{�ï����*�h1�J�ɞ�c����	�v��s�'�E��-�h�B�gR���L��~I6�$<��U�ĩ��Fi�v�k֒���z�x$�W��l��˝y^��K+T��CNx���V�*V��nFby�Ԉ�bG���3i�u��cc0�.gXKށ*= +�v#�P�j� ��y�J3�������H�K /��'�ل9:m�EM�AɊ�v�5O.�Ƞ������]�!�a�FD]�g�T�8;�LQdX������n�����|�H�x�
f��q�bs��^�N�)�%�����[bR��ڎ��h�U���w�*W�Lz$B����ߐAۙT�W��u�s��C{���X~}E��^�%�X'�������w���7�w�,}�\xz	�Q-���E.��4�s�n�F|��@KV����fZ�J��/'���U44�Ϗ^ ��q����縺�o�{�<�:`��I���'14n;�<�Q�b$�L���B�&��w�����'��Ӻ���hX���a�~z	�D*�a1"�e2Իu'�7���;����<PSw��D��R�������)�ڏ.��OYWݶ
���*$��W��W4�F�Bwv�Wg��.ڛ�I�tmM���?�Q����jpq1(�sw���앣��㩿�;tq��+2��l��!N֤��eOsI����h4q3����Nt�����~S��f�{�� V��i�-��5�	�딤B�c5�Ӣ�z0,鏰�lG��l�ep B�|%�y,�UBJ���B�v��O�y�SU8�NK�+���[:k��T�H�I��b�`�d�??�9	�ȇ�~��u���eTxW����/di�S�^"}`�UDc��B�����/+a�q*F���7������?%}�9^�|��D���mju���v�g,{� �q5�w����C#��%|,?���-䒲�Y�_��N�1cZ�~���'M� �1L��7����N}:�>E�B1����v�<1G�}�pz�{�b�\��yq5a{E�R������J"���>_�y�D<�w"�[���dN�*��Ȧx��+�S��x���S��ښ8ȡ7k=�r.�7��Z-�������륑�$��[�_��6�Z��g�����e�Y�To�m$�}]���A5������ro�<�Ue�Ha�9���F�O�1F	��ƌ
����)1���A[�o�&bD^1@Ȱ�TΆ�&u	3|�/�,��`��b��4e��J��_OUV�~�G���+����|�fnu�^�f�T��GU����_ݥ^%��l�T���T`L�3O��kP�j�B1��a��FG�OD
wȀ�Gk��Zej��RV��L������w�I�ehȰ����l�d�L����.vh1=��J�͑}a���|��OU��#7��ٹܱ���'�3\��4Q�ڎe�%"�/��I���·A ��2.�����6x����5pҕ���������s�-��w�]ߜxӗh�T���O$���b�{�z� ���\d�y��?	�"�Z�'S'��>i�AT��:��Ҽ�_����"��l�|`���
������п���+.�RQ�Փd�E`�7�a��B�J�����!W[�<��=!��lw��y�7H��i5�� ���>������6�k&���lOB٦�wHvf1��N�A���&g�&�;.i��E��}W[.�.�D;�ޣ(�ن�𞎃�)�3ࣟs��#`}��$+��K��_��.�
l������g�_�>�%S�NI���Y�/n�&��������Y?�Y���ݗ��v�l�����Ȯ<$�� ]ՄYI�e��d������i��;*O�9�M����-���Jj���Bx�3|#���b���ޕ㖯�ڊ�E��6$x��4����B�ތ\�Î��O��r��c���spʫ�M�q���M����U](�k��&��H��˕V[�XԢ�f���Ju�����e��e,���"$醧��!��lx��:�~�R��A�V�ouSzs�l3�&�BG"U�hVu&�1�h]��!�=��B�鞚&����ɳl��t�E;h8D�ř����C��@ںcL�礹���ػ�~8D�N��gtm��dRC?.�Y�u7���L�9f����F��Mdhh�|��<*���n�/{��@$�y{TR���=%��L��#L���!�툪�W��&���5���#�j1?�W��W��V�属��6�`�q�4ݧ$�WG��4D���[�^%��]4@5u�͘"��O�A�3b d�I\+�L�9t�k'&.W�є~�~�ftT_Y�t��gm��ꄓ�W�4�%���f)�ե��ߙ�%6� �����W<���&H�Hu���A�CX�܈�{A8�!�Q�Ӌl����q�lXW�vuʖP�ap�xw�N��PIDH�|b�6�2�"����N��+��ݶ(<�c�{ Y�`����yr�,�N��0���%�x���}�������E����Nd)t~;!�s�,.SV�W1�T�،�.�����ƃ#n@�\7s=�W�4�����U�����h΋	��	DBdv��n9WAJ��@�;[0�9�>fU�ళ���)�[���Tm[��{�g���V0�K�s�$��mq[E���" �+����2�!�ɀ,�o����V̝,�Ʌ-ۛ\���F5	^�5TK�ڟx�3�5f���X-�t}��/�M]�l�m��~�?��Ɲa&�<+K)T��U��3+�l$9������������Gޝ2����+8�骟[�}�k���=�ZTX�[Z�+A�ަ%��?����ވ����>��m�J�ii`8{)=���
���� ��;nCMb�m�����2h/}��gd)H�Gv�|O�(��γV�+��i��
}+S�!wCa���C���͏��RS��$�^�����V��������j�ߥ)���w��W��Eه[�?���Qr�P�lM�ｹ�1�Kt��h�MR�L���Lg)c�|��`)ˀ��1�7���N��e�,xo;��x���c����oA�4���v{j�mlY��v�����E���&+4�2�_�UU���E��n(Ry�5��,<	�J ��>�����eY(X��8ƒ��8�� ��߯�l<_^4�h�N3A�6#oٮ��!����陴���1��|9N\@�����dK�L�<^��ӗ��H�XEU���?��AXH��V!��K�T;��S	p`�+��*-�M������j@����)��X"���t:�ww�4��ʻ&*�É�O[�j^�o���.���K�9,��J:������[t���P\r�/_�)��k�����C��::��b�5�� ��1O��ebl�����U.�G��kyժ7�� 9G[�tٞ���?��3��՚���-�8O�O���&��Ea�?
N��旍LE��%�}ܥ��hV�����`|���n-����!�%�w8!=
#z37C��'J�2�b�,��#&�zFZQV�W��~tL�򴒟�kݻ�ޥ��{>I�*qk�%�9e�%�u�#?U{z{X�:�	_bty�4OA?���-�	�~
.:+�C�c����Y;��ݭ���"k4���/��4mO����Aza�4âI��X�?�'���帷��^7r�_���?�L/�4N�^ʌ�` ֧̚@�����}�Tl��Tq"氓���,Ek5�H���C)�������T _���0P0}4�25��r�s7u���W)I<-vN�\�eS�fzh��뢺g?���Ȇ�d�H�%~㷳���	�~<��~�1 lY��b��"���R�p"fv��o�ןQ��sG�T�1p�%J7Dw�_����÷��y����B~��NL8N����R���岡v�\.���\��O��n��L���h�r9�,����=/&���J�J�fZ�m��΀q�傎���$�R���ϒ.�v�U���ﳩ�J_r��8�ɓ�b{7��,���LY8���lsQ��3�� 	Zw\����*TǯU=�֦��7��d���٭��:�5�a���aZ��.ׅ}"��D?<\�ɟ󊸉�˒	�ZGp+غ�o��wjo[��:��BU?(����X`]�L ��X�G%ߣ��ꪽ��݂^��X��:I�㧚u�~+7Z�(f&v�� ~��WS�t`3ks��ő�ހQ���t�5|:���:�btm���T	�V����u	������b�@^���y�� �z��{d���iNy��"����iL�W!�?\���}@��&�wō3%�W]w>������M�_#n}*O�lf�ıvp���ݱ�q	�f�*S���������(�A���	�Nx7��;:^_'�6W9'�9�L�3��=(|=q)���$�
�45"h���7oE^qƔ=��o9�i���@(����A��P�������G�W���X��ƪ��VG`Ƽ�.�������uٙ,j�}�/�e�&j.:~+Vw��Z�8N8LϏ*O6g>�Cs�W�U��N�A�F03�"�,b~�aH������zA��%ɒ�����L@� R��_��B�җ�
�T�?�<�$_ʎ�(���,����*��F�PU$����j3 �DE�ެ-�B���2�,?���G-�1B<$t��6�:��j`\v������u�z{z"��;�F+S}`m>����[=�����H��b;�v{N)��}I(L?ߜ��̉֐�t�8靤���S�D{��f4o���m[8�/l�W�T������M!����KP���\�a�*eo��_4�4�S��3��{�A]�0����af>ڇ�B\�M�Oy�,x��d��i7�:�#-��@_��X�j�N�`ב.���%�?�;K��^��6�^]�=s3p��l�� *�|��p���6���E^�xJ9ct��0��^)@ʪФ`bgSB�l��t���fK��^��Y��q�!@ď�����H����~�;QI��2΅��>��6cK@Eף]G���0bSofo��Ы����(��D��j���'�ѕǭ#�~O��_��|T��ՕiiI�Ȗ���w�d��=��ޞ�e�g������wѹՑ2�)��&���`���	ư�����˼��"��wO�Ut���&�8Ol�4�g���Z���(�J��i� �@��Y`}�Q�g��$�������y@�����t|��ٷ�)G1�@g:$�	�A?�)?E�zP<I�<��5��(E�-���e�:����g��4�؀Y�S79/�6�v4�|�VR{t�J]�3c4j��&o�>"	�F�w�e	�QfE�C�cx��w8z�{���@�b��,�:�<����G����P�d��C�����K�}�����Rxߋb(���8fo#�N��B�h?�uɍ������ �
��G��cl�#?�e���4��,1���q�u��߸Bd�L�IҙY��cq�)��&tN��znT��L��GN����͠P�O���u��
F$�Un���$WV�t�k�,t�d������y��=,$7�v�"�A���S�ĭ���+��n>�7+�&�n��� ���oL⦝.�&�ND��q!Y�D_iQ׮�S;�U����ɘelO���P���N�Ic���E�}8L"-n~eݪUg�K�,���vp�h��{	w��?���|���l�����z7z���9Ȕ*��c���hi_ՠڌ�QZ?�@i;.��kv�4+$�q>So��+�f����򢥒���b��o��><5�9�����.��l�_׏s'�r��k��)՚�S���3�Q���.}v��j�ݪ&{®L��=�O����yZ�L)1<p����p�ĭ��y�c���/��c)*(��w|�s�`�?��\��3ل*� �2��&e�h9w���ɫJ��*��?�Q��D��V�W����mi��<��)��^�TK�a�/��=w�h6m��=�9��l�����B��GZi�Xi�X��ɇ*�M�����<(n��TɎ��S�Y��sC�1mI�d����.���t�_�çJ�~��7?L�����s���E3�jJ�ǌ��w_eH���ϋЇ�-�Z,w�d�<���q�[��_�^�P̫7��~���XQP`����{��#:Z�sZx�T�;��źC}oߗ�-C�fS�s�E�c�R����[������[
�rqߟ	O_��V����	>vʮY�_�`�`=�G_�IS�Wmh� �ߛ�;��@�s�ݕͨ!i����7����8�+^�x�?��V�����/��b�,�Oq/�q�8��a;�ZEɱ�H��Y����y[�r��D�~6���ο[��U���~�̋t���9�i�w|�X�3j�3:�;�5���*(��9z� �.�菣����*���V�$%�:A@7��b�T�/M\=Q�4y(���R���!J� T��ݽ\]%�hh��-	�9t��>��IY�j��APϟ�nSo@���\�D���e��������1�8q!�50;��J��T�4��D�$�QA;}:Z���j�&�x��l��>�f+�v=).�i����뼦n|*n��v��;Ƌ���1t{Y&�P$�O�5�&��"��b�a�v3)А;��.��UMȴu��ih�{Y�v�AuA_��K�Q���j|�	�| �iZ��YK��"��%$�q�ߠ^YeR�`&T�oQ��DH�cv�g��`'���	\9�D����A854�~�&�Y	<��Hq�iR��W���]:9�����+V���'��7����>joP+k������>��d�e��N�!�����XGܛ;�#�{�l
[��u�8���prr�rǪ�+�Y�|�T<+W��@���ǅ}62�-t��Хy��&�Tʭ����.�&5�&U(�{+�^+kSACC[��D3��}X![�E�{Q܌�V�.0�l�ص�5�˺K�~�}��m[ݙ�Z�F���y���p?ջ�Fkx��-��9��_���m�[��ʒh�`�v���7�X��s4��Q��\� }F�d��1
Y,��I;�75=���j�1m����1/?�� 8�Ҙ�2�}>M�R�̽]-��������k����c�Mn��Md}W���iul�	-�)[@�[�BV�G=�>�rB�������g&��U��S������J%c#z�I����͓jp�w�f��-��\������v�Q�?�-�m�]��<�!?�%W��h*�s��;��a���GN��&[���]��@���� i�����\"��.�iTT3�G"���D+/Mڴ��k�.)w�]��d��.�0tZ��q����l���Xu��1��-��',Y�*j�:�yT~�j��8 ewV6�c�T���"�	����@���M"��ܸ�P*��堏wj֙���]mV�X��쨔��jXM}��C�7�����c_��b�.�2}�:@2��f_lq��/�:��/E~�N�FX��+S$b1Y ��M��ξO��d��bu~T�I��J~�_[�l����@��ݳs:Is�#@�h*q���P�:��而:`U2f�I��U|5�{W�����l�	 �7$�J��`�r���.�v���'D��4-/��G9��})�Ɂ�{;�u�Z����(����q0|�׍�zm��Bm�Coc&`YM#_��E���{`n�^�W��*��4�e��}:���(���mS�1<���8)߲�e�a�G�鼉lw�V��VA���iy��-������e��^o*V�����U�^��[o�>�a�I��2ީ�Љ��¤=���c��.=��X�pe5�݂��u��Cz�ڳ�Җ��8�E[i	�$���Fݼ�O��� g{�f�0W��#ԣ�j���"8*_7���P�-ձ���c�(n�ҽx��H��t���NI�K�Z���2��e^�e0�͟�g8hh&���8�R�)�� ��J�ㇴ�K�k̤gtX��X(�WC,�r�n��G;3�ot<��o�ʋ��@h�u�DO���o�x�鳧鲧�8���zT���\���.*MI�ѺO�Wb�h�a>�1=p ��<1����:��$�-*�i�S������fij �ۜ�;L�z�<.tc��O�@���x�?��#<�����$���γ�:�V��J
������PK   �n~X?�]��  z�  /   images/0769869c-6d33-46eb-8102-928d675c2604.png i@���PNG

   IHDR  Y   p   �&�   sRGB ���   gAMA  ���a   	pHYs  �  �(J�  �IDATx^����Uu7�;}�ҫ��t,QR�c�1�H4jꗨXkb�%�1F�^���`A �.l�ݝ���}��>����l�e��=�[�=��-��vM��-]]]���w�n)���=������t'�Iw,j3��&��9Ԟ���g�67�ۓn����(6������U� ���2��:�m��2����j�{m�͕��ʥ=��u3m�^:z��Qۧ������r�9��
����]v٥�����kז���
�===�9�U�ӳMvo488X�Ν[����jc!��%�oid7�sNF+V�(s�̩��d����Z�xqձU�V��vک��>eѢEG{
w��7�����_��2�sD����������H�������~t�N�}(ےn���կ~um��m���:U�}�ӞV����֊̅��������a�K`�#���$y`�p�{޳��� YV���_����v�ae```�n��#cl�t�!�L�u��K��e˖��+W���C"7��k��jǥ��i5�D���볽Y��Դԛ����G<b��I������E���O/\p��e["�	/�#�<����������D7~����>��5�4�i�I��m��<��u�YS�]��F*�>�Y�*�������^�O�c � $�/�59�y��HyN=������S�\����������������G=�Qe޼y�~IK] ��;�\��ַ�7��a%�����U�(æ� ��ӟ�ty��_���~�: %˔�c� �x�;�{��[u��NY������mo{[�ԧ>Uۧ���[���ٽ��(����˃��r�WV﷝��|�ӟ^�6}y�s�Sv�m��������w����~5��U�wJ������(_����v��#Q�SN9�|��_�C�T@I����r�W���P
9��mA:�s�=�|�;ߩ�	F�$�caX�WϨ��_������-����=5�G]]-����s�I'Ն������~�������O��O呏|dy�P�+#���O~R������z?�'P�7���U��~��;���D�'�@v��?�i�������O~r� �+�GuT���j!i%i����w��xFyғ�TeKǍ&:���'�\����i�e�n�^��t��f�zha��Bg��l�m�j�)��-_���kH��Y���
%�@���rg��6�[9��h�r6yɒ%�[n)���ãexd��^3T�-_Y��tK�ii�]O�-�,��4�+�^[z�j��u2�_}��ʍ7�X�^u:7.������W�&�KwoO=WV�5�\S.���Ox�)��	�)[J�=2���4;�����6���H/�K���-�_�GGJO_t��]e`n���ͭg3�dm7:6q+n���7��n�{����v���$�÷�8H[Uq�l�{M��PY ���	��xb�Qh�)s*9Em�'�潭ɹ���FF��]���%���?<�04�^'���n����H��kH�G�-(�cCe����`�@�7gn�;0/ b�@6���y�?�L�[�֎���Ξ5��4���=�Q�7�5��j�������s&&�$2?�~�/?���g�{l��=�q�O��2�}kY98T�zB)�ˮ;�Rp���S��g�O����'�iyʟ?���.w	Cn������k�m�y��m��ȹ�=7�d���m�i��0�~Ɵ�3�����{�3�YG�Fm��^��W�Q�鹇<�!5��Vd|m�N��m�4���y۽�Ǚ*�a�&�����D��p���j��2���ee�����`�s��S�lc���`�ny�Cɫה��#�VW�;����2��U+���PY�|iY���2l�dh��\[�#��{zB.cy!�H��^��]��k'���	R�^صg�Sɝ����A���M�����5�s�9�$��<{��fc|׻�U�����͑��Dȸ�lwY�pQ�ǿny�;�Q���o-�|�[j�g<�o���jN�t��R<���7�����//�|�k��_���ʗ�{yȃmo�e��^m�$�NʷYܵ���+���ްS2��@����^�7:v$FtCC<F���2��8�e�,���kc8ә?a �����S���;�}�f	�
}�_<��r�/*���̰��ш���vjם;
՚0&F���u�]�����[EiI�*�|�5I��d�p��0��������xKy�;�R>���G?��2'<X�n�I��%;������|��-~_���(�:��r�M��}�F���b�9���{��{�V>�_oy]y�;�\>��w��{t�2E���]:��|v�����>�|���s����+ ����ډ����ʗ�ɤl����+��	�Y���*������s�2�M�v�{{�w9�Ꜹ��[�8∺;��Y��e�nMY�zY\v}Y����Kʲ�/����?F{��>Nt���6:��5ˣ����tu��eͲ��ڕ7�����1B��F�*����r��x4� �s�F��q�S�Fx��C$G#3��Lz�5���f;#מ͆�#����:�ʸ�{�=�أ�aN���'>�Ο7G��U�%hB�<�l�fe��J�+��z�ƴ`n_y��ǕG=���Q'?�<:�Ox���A��YF��������+;-�_�ȓ�c����'�\~�C�^���<	�
PE����6Vv�iay�cV���c�����=��}�(=e��a���8��:-@a��2ٮ�����h1��R�6Dڤiڬi ��U��8���Zݎ;����2\3�͡�4����,��5t_X�3����~��4V/-k�_^V-�]�����_V^����׽"@v8�8�9�W����˚[�,�n���\rQ=�Y��L���1�GۛzB������+�Q;�'��c 爄u�a"CS,M��a�%�m�����~9f�ӑ�N'y���w*]���X�~�����%����������*��e �^15���7�#S��cO	 �/7\yIYrex1W��,�����.(�,�����014⡄��-+oYZ���/�3���r�׿P���ϗs~�ݲj�-e��9գi�:�ԣC�����\�럕�.��\��s�5�;�,����p�l�S���2�����6�uU�����+���P�!͖Ի]�q�V�Q��i8�dXƇ��򹰌8��~��%I9LUx)���t�</�*�p㣥�'�0:����+��{��ҳ��һvI�^��t`���8��p:���2��2>�������.)c������#��m��*�X"�m�}�\�q�0�|��k�S_�F�Q��tċU��<�15����w߽>��n���¹1/�mu |�k�퉪Fi(WQh
ӑ��o/ja��� ��{�0��W.-�+�hV�P�W^_���w�,/szM�x�1��Ck�՗]X������/������ee{C %vb�����)C�n)Cnd��f^_n�f����5Z�ՌcO�6'���UW]U����o}�nW����/�ŬI[0��f�d{��$8b�V[;g`��=-��ܧ�Q�cq.�fڛC�7ѻ��H�<h�����D?{F��@��ܨ�������Y�j� �hľ�̔�����K����71Tz�u��d�:���Mٴ����Җ�|�o�7�RgE����zx��6H9�/�c�_�l'�"�dJ xJ���&�3g �ym���-��Fy��|�d*�UM"@�dS�����|{���qt��Jo m���=�����MoO��P[(`�9��pg��zx�P �`�z4���p�Ll��U�$ؚ�
��vM�+�#npƭa[�� �5H[������f[;eۡ<ϸ߰�S��g��q�3F�4�-M��$F��U�ɮ�J���x�b���)�'<Ѐ��I�S�N�3�/z�������@�hGK_����/v�R{+�ݖ"�@���v�G�V�icm�S0������J?�C�d���N]�� w�ѱx�Z줚NQNQ"e�ި��&��4��H�NX�����R�g��:��5�l�G8T�'@6�1Ƙ���1T��3�MA��E�C��u�a��h�ue��S)<��h=�h�ed<8��$��l3��x�X�>C��i",=�5�!<��g鼙�lmsH��{8뜆���Z�LƉ���M�/kcD1�?�_#\��7����hw2
}0�`q�+:�VG��3��)˙2d䢝 �s�ia	�
�Ӥ^6���a��<�C»���p�_�g"qs4����). ΰ��퍪֦����h
i[%^*`l*@K�Z�P'
Eq�WЉ8���a��	�����BV�nn}L.-COb�-rϬ�M��n,e�<f������[��}מ1B`�(��n7�tS|���,�^z�.r��܉����&պD��{���S�����-c}��hϼ2��_���=V9(k�D�)���f| @xN��+#��c��UO�\"h���V� �$e;�]�k�Y� ���Ԧ���8w_�:O���H�=�m���f"������s�����f=��u@^��ިV��㎛�<��7)���9T��YD(Z�2�]1,	�u�kN
�ꋚ�P�0HyF�\I���0̉ed,�&�KOi	C[�v�z��N�,�u�x>��N��I<q>�s��'�!JEݐ�v"F�S�y̶�g��s��ò\����g�YB1u��Б0>��)˪Λ��g�ܣ!G����輲b�@�yeY1<�/,���p��J�u�]]!�h����s,+{�*+ˎeu�6S�@������C��N|{9���7�h����f	�¸��sΛ.O��6����e�&�ϖ�������~)����(]����^YoZz�R8e����FM�_����{�4ȶK-�1�� ���6<��2����1oQx8�=��N cx2��1�,�����������kBQǺʜ��k�&	�]����{*�w����o���x ndTt�D	uh�{c���7��y�a�L�� L ��P��<����T���c��8Q�p'r_y~r��בN����+{�{P���{���=��}�{���{�#�ݢ�dō�e��20wQ�y�C��-�����~GD��C'��}�xx\�1ϷEJ�hmb�5���������щsm���di��8GҕF�VK�-��+_�C��K���`#�����\z�����}X;Pn����@U���j6~�<��}Ki�[� Y5�I��u�k��h�.^<���y��?�Y�pvl#,�����XwG{b�< �??�1L�:�DWE�z��Hs�ҿp�2w�^e�N��w���ۚ^��X<�i0+�:1�o��# �Jh�s���~-�Lo1J启���V���9WV ���4�<�\n'�J��Y9Qm�`���v�a��h�}���R�_��>e�=�o��b�E�`o4y�y� ���{�2w�Ne�]�.;�W�u�}B���"�6����9����h	��;jO��&<�sы�CR��!�(�9��~�H��k_���A'����E]T=[o?J_�|�n�7�5bp>��A����>U�h:�j���zKP6t;U/�N�G��� ��>��w�=+�{�=˼�;��y�Tᵎ*��v��y�s��>���3�����9���r�!GTOw=�����C�y��Ï�y��!e�=(����Q����+u�ϣ����^ٯ�����F����W{�{��^��fO���4� i3�<�4��b)3ϕ�Qj��)��	+-�,�sq�I�6�ls9)u);9��Y�X'�5��[n�yY���>Y^��ה{�k˿�����������J��d�������U�9����W��<��//|��˷�����{��ڦ�R���>�%i_���-[d+|�D�qޣG�KMJ�	瘔�g"���x�/x��W��"��	�2m���}��Jm�Nl(�;u����j�U��C�M"��|��pzL�=^;b���u$�de�.�k��f�֎���oZ��\{��r]W�
���e<�si��,*�]uM���˯��\}��ep�������F��$Ny������%7�����\}�-e�M��uK������W=Wa�j����=��y+r�j����#We74�ͽ4,2�Q`�p+���2!唦g�?���u�AniWe�rgz���?�q��?��[�!�r�^5X�+�)�o�yV9�?]>󥯔O~���+�?�G!���oZ:����'��|��_.�>���g�Y>��O��.��,X�x=/6��2���7���Ѿd��+�qT_:�v�ژ�\�#ap�7u�1۽:_<ay����җ���v�iu�s�V�{���=��� o3�텺Ө(��8��!� ��b�)x�0���r����c�9�z��P if�v8�9�?��r�'��Փ�w&j�fw��k�����?����'�ey�?�<�я/_��*ׅ
�o�藿:���S�V�����O������VY�rE\������\|�e��O����'E��?���S��<��O.����
�����������l��'<�<��O���"��vKb ���e��3|���5�8��xiX���@~�1bm��$] ���E����u��y۽��e���[ʡ<kT����܅1\^�CY�h�2w��[�t������u�}��Ee���q�O�>��Ȏ��е����uu%�0�%3��B�[�l{�MN�to6$|��N*����������Ճ�.��>Ϻ(�t�qG�@��X�g0��?��H`����WC�"�0|����<�I���q�0��CՎM�ʩoN6�~�k g+V�.+���W�-��$o^��,��S�§!��uY���[*P���&��(k S�� A9&�;�e��X����e4�a�Me���n�����6KL��I=���v��Ɛ�hY�d����
18�X��#��gH�LC�f8G�\<���I��hHz�9��EV��ENi|���=���Z��b���$��%K�������D4�CT}��HY��]Y�rmW�Uq��m�����n>�Ie��l���P���͕ñi��vF�	�y��qS됺���s8�H��Ka��ݞ�kbtlbe���W^Y�p|��m�x{5LHC���a5����D�RIK:fZ>]�'Y|�<�و��}���_�B-��!���C�s�._���+b�1��
n�4�P(�y�s�Ñ�����G�o[y������=������0�׾���ǟXN8��k,����)����5���2w�/:#�Bl���e����y�Ax�O)'�t┢�����[�l�!y���B�Ƅ�}��Qh&j�2H�=r�=��\�<	�x�ڏZx3Vr��ʼ\#�w��]�1g{l*I���WT��1��k�_���O��N�/a���������[sx��E�xB��/{Y�e|�w�ޓ���pt�~�vd|�~�������������'M75��UuiR>k�A�p�?�0eZ�g�wO�]�x�:��~墡g��N�|���D�xtW~y_�8���m,IGY�|tV~�=���[��n�I'�H ;:�.(������]��9n�J��d���o���#�ը����B05��G�t2�|M/�w͆wN1��{�>���VOld�5Y?���+��\?�x����&� ��a'?"���?�~/�7��u��7�Y�c�J3����S���޺H���0�� ���7� P���5KV>����O]k��g�uȣ��w��Lx�V[�\�|ս��R��K/�*��1�ɇ��O^���s�=�6r��4��c~�x��3�=K O���K9�����l���k�2�d]y���җU9~���_xRm�ìe���-��XN}���P?MϼV��qi;@+�7�����|���u�"f"�����P}�~��睨S\�\ۑ;h� 2,�%�#�֤��NϷo9>���)oS.w��xɋ^T>�ϔ����h(��������v�>��w�c(���o��eXGS
�r}��q�lpi;�������/���{Պ�Uu^�/x^M��!�ׅ&r�-������գ�����`}���<}��9�����r�ΙRjsį��Z�M�6L�Q�$x�_��7��+G�M�țq�����t[^�9�W��U��u�hډ��2���I��t8d�)$Nr^o��}L���C���ՒP'��B�NYG�~r楜�ӏ[j?�����z��k�id�1��ܯV��y��-�D�R��_�E�1ډR���c�1ډ�=�sA^���W5"�vJ�6%+ݬW-O�i�g��!�Gc2���s�K��>��r7�ݤ���ٶB��NU|�k_�jeN�ޑ�z��e�K�W_{M�i�-Q��d�ߪ�x<,T���ޙ�v�	ÞO_���@OSRyy�����\�`��C$<J�@�W��*o�����)ڪՃu>���	]#8f�u�T���=�{�h�Q:�5N/A]��]01�e��Ԇ�º��xމ2� �,��k����C~5�F>�r�0d���k����-�7���3t�shڊ��4,����~��W;+�:�������`���=Q�,W�3�($S�o}��Ѧ��Ԭ�a�zbr���}�t$��^�2l�i������|�2w����9'�����g>]�N\���F±G�[r�u~�<�UZ�xa��^欩;J��Ѩ��e�\R�����K.�?M}�5� �b/y�K��$���d�tPm�s�9�����ޕW�SA�������g6�j���W�w�g�t��=�W��僡J�j�-<-ѷ��4��m�������� XCW_ߨy�����0��# ���y�w(�#�<
'M�\�}CGi����6�*W�K��φrS9@���:`u�[MA���?ֹxe�>Y�$q��o��o�>�L?���S���G��2ފ&G(��UY��Ԕ�4�>���6A�����ʑa3�k�;ɵ�n�i���ȑ��	�fD�金�=����0ڝ�4;����o�m�;�:������O�R�m��3|(��u�r�!�}������hQ| ���;�/��y���R�9�W��"�s@A)�c����0�^X�<)pS�L�y>I��I��Ґo�c��ř~������˿ԡ��ª���/}�Ku��px�7o�ze�_DPGy���)�f����,k�ڹ4���EX ���m��I��3Q�e����g�M����&5��\Z���ӕ�模^O�K�l,g:�ȓv�����4]9;Q�u�L�ڎ�q�'���/ =�������	Y���#�ډnǑ��9uGW�XY����z]G��F��g/�ێ�)WY��9�+|���a��n*>0�F@�q���N�Gcz�����M%^XFk~�0RZ�I:�ca�#t$���8&7��OG�\��W~�L�yД�RS��_彫;�S�)�t<KCPi�?�P�@	`XG�e��IY���<3��6toK���i2Rm쾲`�7��������g*��[�7����&���m���v�k�s��f��~k���f9g���u��z����~�nmR>#Q#Y#ЙX�,N�	��EҦ�ѶF]�}�Z! ��o|�[�MozS���<��

<%+�3�ɺ6�7���(I��]/3H�6W)�{~D�7Ș��-N^�K��#s�3Q��&��1�ڪu=F�Z�Z^�{���r*L�;�:��幸�␁#�8R�3���s �Z<�od�C �������0��=��	jG�~��^Vu��ޔ��G;Y���a寣�Ї>T������T�����)�@3M���.�T��P�ice�N��PvF�ֹlc{��]�^E7 ��m��-�1���-G�.!�;[�����P;��(���p�����#�y�r�_�e�V���NU���dR��R�'�-A�qe��-�P�4l�arO##[����֕w�!�|�#되" ���(��@ @�ꀳF zfF+�j����5����e���*�����d�ri���p�/��qN�<Na3��W�k� +,"�!�2����,+%u�Y����?�I�S[�V4u��H�;����z�݋�NyO9կI�N���GV;�ӆ�x7���9k_�⩒3�Ie���yr�l%G4�`�ͷ��o\Z���y�,C�.+#+��n�CY4����ZC�k6���sW<���3������D�[R���7��#7�9#�J����=6X&����xY��:����7ڻv��ܡs�%��ň��['3�rp^{�|޸����Y��0Ώ�g���(㯣��L	�Ƴ���c�j7��~���s�� � `�a�O��T�jNҴ � ��$�,~�<	\Z��Z���x.Mf�q�m��t�ʼ����8I�=��P��1�˱~��-�('Y���X<!��3&;���d��$>��4.� G��ܟ-gY�/� xZ�{�_��W��w�;�/�Y� �jk#��7��Y甭����'zhzS�ȣ����S���Ϫ^�S�򔪣v*,�����Z~��s˃�9��U�|��k<����<z���4�NYf�Ԕe�u�K"#7��HYنrsF�M��J;e�$���-s�P������k�S&n�Q���3��{�R߷T>l�Np���q?��>�x�R�9���K��9��Z���o(K����3��Ug��r�����ߔޡ�KO�l�Dˆ{��UCI��1���j�/�Mr%uzCqkE�%���MU�
��j����2�ֽHg$@����~��L���ֆn�������|u<Sظ���ɉqQ�[�5662���m8��PoxCk� 	 ����ޞٜM�\�������m�DR'Ų׏qJ��g��%}��,.	P�ڕ�V���RZ'�N�x��nM��@������Q�m?22`L�M�	`<sϵ�W��޹�9`$.vI{����N���wl;�E?��E�aϖ�\�kgC�w��ݵΩ�hv>�8SQe�Zy���P���H��?6�?�����lHm�+���G��Y��(���4������P�,�I�p�q��j_�'G�f'�c"���am��.����9lg"�bA�`�^].�������/sBc�������2��<AeMn�nܫ�e�L��+�_�e�����c�(܇z$_z8�fm
�]��/=�e�{n@�@9�ȓ�>�?��]t��h�����g�V�Y]�<�>匯�.xf�ԧ>e��)\od�ځ#���Z�� ��rC�����v=�,X\&���%Kn(��{�����\s��e�?�F_��s�n~Aw��5��~����aw/~nb�-������r}�ļ�x������]Y<�~�JȲg������xr�5�3Oc��#�Hh�!
�5�E1��	e�I h����M%�L�0 �*�Io�
����@Ĝ.�N��Iʹ:��L��IӁh�ƀ,N�L������s�5���a��$�Dn:BL���I��l�	n)g�!O@g���0�� ���f��g�RMY�h����a�@�������9�4�#;��6����g�lm����I�j�'�Q�s�a���4���*�p�u�e�������L �������}�₏���K˼�=e����tv�i�r��M�E�ܯד��~�	x�� ��g�حELD9&Fyy�^g�Q��|K֣�ue�u���˟]�h�}�y~Y1��z�?-����{`�����Oy���T��jg�9����)哟�ĺ��[N��K��nI����Ug�ߞ{v�ޯ򐇕rӯ����n��'���߽_������������_�����R��������)�[�娣���_T~v�y�!�}\)s���_����r�cS�ٟ��g�^G��|l�����9��F����Z�[A�p�~4��}�8)���(��f�VMTSNssi�.��hHúG���$A�\�7���^'jO��6d�+���׿q�igڒ ����_���b{�5�r)����j� s���#G�����.P6���6$���Դ+�^Q�0��4��9$my ��^���f�{�_���7F��J�s���9�S���~��&�}$��o�������x�AO��xʃ�me�<��㘜$\�e?�1*�5	��@�,`�/�Lx��!��1<��e�k~��h��¡-�ݵ��Qw��Z���Z��cU\��\��ؕ׭�p�p���8�s����K�OM�t�p������˚>8�Cx�)�prY�ˡ���|y�[�UV�#�X��g��W+�~�S�Ss��GwZ�_�DOn,+~��r��,]�����O0�����T;6����ʷ���r�=��Zd[��r�����ed�D������ڛ˽�?��^���󓟗�?��w��u�^�O�#sR)k�5�/-?�ٕ�)�85��p���Rcr���561<�W�G�+�Ͷ��u��7��%(��P�v�FR*I�t\�L/
y^�=(�5�ӽ&m,�F�{���zֳ'�v��٤����cy���^_!WFP}Ӷ�ȀVY�2�ʽU|F��O|�~��3�2 �γ�P�!]q���|�(}���mG�f�(ۮ��I	�T��#?���Cx�H+�6��P�|!%˸�ZJ,��1� Yq�<��P����u��?�AS�M�v"Se��/~�T^�Ͳe���3L��ūWz�������3���˷��-��	d������k/|_]}a���ܲ׾{��v݃��©,^�*�(�� �u��0��cX�k<� lJJ�Z�
5^�	���b����������e受��N*B��Pv���rԱ+�G���/�}ċNp�8��{�����~U?�(N��z�:�jM^� �Ľ+.��|�>��n(����rԑG�=�ZT~��ߖ�[Yp�����C�ܟ�_V�ݥ�ɟ�IZsq�ů~Y���>�^�ݫ��sʒk��?��۞�W��]Yr��r�c��:����O�=r����O~|Q��-�D�/�rE]ó��+��x-_٫�����w[�|e}ؤTtGLA1eIr?*�-��#��0�L�f�vʰ��Ƃ�2+/0������|ڙ�4�:�y�^!���'C�%/91���N���W,/o~ӛ�.��#��N�ZPyԣU�3���I:J�`�mu	Ħs,>~�;ߩ޶7���x��= �+s���	�o�p��w��]�C/<9�+�|ͯ��ph�4;�k�=Y�	�=�-	���ei�-����?���?���C�-g~��	Ozb�W�ɝ��\x�QOeR7�$��υf��$�/�����s�����9=����Q��ߕK�}SY}�/��ݿ���ꏊ�rB�
��!,� �+�6@��iܯ�c�qi$ �8q���c���s��1l�&�z���+V��o-�\׽]e��\�st �@OY;�2t:tpde�=T�9��"�Ȼ�.Vp�%�:݉(OXnܛ(���e�_U�;��%+����c ߁��C�Z~�����W�X�������\[V,﫻�֌\]�;���ߢr�Q*����r�7��~���~��/�c�����B�ڋ�Λ�]�s����n��\���~��=�D��2<~M�����D���^xdtAѢ��y�AZ	�D�q&�"0r7�I-Ah��)/�/���mI��~*�&�*L���b_z�<T��sw ��.&o��{�@�$	��׮�/3J�c9���zUyU���׼�5���)��R��Җ�vt����1Ea��ܼ���m?��&�(���	қ��@��H�#�(
pxu��l��P�1��]��?Ӑ>Y��܁�w�4Yx� S�x��]�N�-��� ����=�F�L���3��w��'���DWY����ݯt/\\VD�C�@+Iu�$�����I�$�����y���GƱk<��~в'��1G��`n�{����Bo���s|l������y�7`��ݑgw�����q���\ƣ��N;�+.>Ce�˜>�������Bs���}0ht���)kW�6�m>�.F��7:�y}�!Ǹ�`^�D<���OO�x��"]�����O��=a{�}�IU�ъ�orگJy�QF����y�lH�Tn�L+��{�����A��uz�NM��b�yO �������(x.@�W�#d��k?q����(�8��l�N�&y4��KSz����������4���⺖�k���N��D���R�:�
�ys(Ӕ/Y-��H9)��['�z��}���i��7�~�NS��/����e��e��pC��秙�|]eǝw-s,p��(v�<��&�z�Y��!�܊&A�29��<˄�����p�; ���;��e���W� �xX׋�}m`���@`�[�u�w=9=xMY�󚁮�[�|ͪ�N��֮#�G���P�����9O�'
pU+���^ 	����5!�(Wo��G=4ב^m��o�ju5��<�!�6Id#N偹sʜys�G������)<e5��MX{�U-�pN�	 MJ�Bʏ6Zl��a�n��/��S��q:&�M��{h9��k��Y��+�}�v�gx,��-
�^4ٞ�E�p�Eo{׻�_z��e�;��q-&�̏��t��#�����yX#.e���x@�鍑m�+T O1��=�U��iW�r��+������e��Y�)+F �42/o���Q'�M�,�����x��NL�ȑt`t���y�z�ʗ����N��W�����pHs�|�����ᑡ�0���ΫAW�����������;��oYV����k_=�|�s�/�������O(Ck��xs��#��tܪP�qo�O�h��{��Y�]vZ�S�����B�IyM�S"�O2�,���|&���G�h��\��X�������v+��Y��Z����8�e�t���L�c�g(C%�%�_׶5����qZ��zx������jϽ���Dߜ �h�o��p�p���]ƣ���%+��B�+`ׅ�Ij�d�#C��3��̎��SO=��_50g��|"����z[F�b�O��������i�W�|�����z2C��K�!rQ �4hrÞe#"�K�	v�L�<��.�oQ;�5����|��⇯`V��r(S�/>���*�7Y�ʙ��2_rwL Dʍ�wI�����Km��4t��F:ʧ��X��=�y�Ql)�ъ)`/�� LS���`� M��g���sz�ʪ܎y.-Gr�v&'r$W�]������홗<����$����@��rO+�c�<lxn~	��O��k����y��j����t=z�֍+�	�玭��:���8��k��)C�� ՚v���;ʰ^;wQ��>�މZ�c�&�(��/�h�z�7�}�?�A܉n���e��[��.�ToB��ґl�&�>�'��w�B�� U��P>�o�8?�m��'@IM�� )�mD�p�V�����tl�0��L�S�=���nX�1���ҫ�bdy���+����ms��*�'�x�1l��-]�*.�"?m�09�t-�p	$���*p}�:;V��������=m�9v?���vrTn�X��KpUeLc��Q]S�~&݋[�������._uq$���o�59_'�o���mE�LL���봧̫�l����䤦��D=1�o�w��ȿ�C���|��$�# l[@W�)��O�����4@G�֕� ��_�IUGk@O���qF�ړ4��oU���אab�"�"��ՋV�FZId'σ�CT���uO�{�z�0ɼ���6��>l*���ܠo�,U��$X$^��-9I�UhAV���J�BR�v��������f����� ��#���(+c�
L�,��g�	�Ƨ�	8�>M�	��+�7哆����e��v��n�䢈t�+m ]�+OX���eb*�waO<�r��V?�n4�WL�X �M�/�.	� �GgG�-eF6V����[�
o[R2���/|a}-V:ꬼ�%=�cu%3�L�l�ɪ�N����K���:�i��3�d<�6�D�#M���.�iOu�6�l�N��8d�d$N�8��Y[���k8`��[I���}�2L���
*�N;�xڤ
F��C��K�*�EgP멜y���ɠIY�)J�Z�SA��Q�ۉ�%&�ԕ����� XM����W���>��R :@ſK)4��0b[�(XzN~�/���;���a6%�p�D��5w+E)�-C6���d�L�=�1�3e��,��AަB3Q6��5�� 
D�/���{�^i�ع� ^�a��a�/ ���Af��2�;U�amFv�N;�
v~@�ܹ���>�������M��*���vU  ����������V���^/zы�^ٗ��e�u��������w�#�8�^;b;W�ɼ�)�O�FV�����	tbk�t�.�/u	��R/��M����''km���:�k���=:)m%���M�  ���i�v��:�l�<6);'�p��C��:�ex�2�v���D�m��.�hhnJ�Rk='��e)Aw�ìi����kTs�/���b����# ��];RJi���f��P>a�j��zoS
��SH�ţ <j@A���6jO��/�� V'�oRI�TNL�KI��]��XȎ2�<w��D�����m�����|k�A� �)��s�^2�_Y��v�Wy����[�^��&@�>]i�\��C0bq���?�n�2갏ֈ ��F���-�;y�y�H�ޛoH�y�7�|`ƻ��2&�\{�S�_u�v���nd��ȵ	������-{1rs����:��n�{���ֶ\��\y�U媫�,s�Zt�UOoY{Jw؍�Ŷ;i�fnw64]:ѱML<��ϫ_�gd�W�Fi�!�� �}ٜ�^�F�Y^�Π��!��C�Д��`�x����(I��d����d�%Ŕ����Z�����յ��?-�7@>�	�<�9 #��WW� �$(��9�t(u���u�d���.`h{CY�S����*@��7��(�CSN��K�<J2 X��'�K��9�VWa�G�Uv�(e����t"��J_�r:�+/ټ�(�K�ɟj�����:�e۹@���,����n��RG���3���l�"C�l����L��,g��E��cuۚI��������l�/#('G*��x8"���hy�I��	G�Sv���i�����ݵ1
��N�q�S��OqG;�P`�D�6�~-�DxI!#�}׀MIx^�y�8y݌W��F���bl���./��V�>���0�ܭ1�儬)�!��ՑO�bM}���zyK/,7t��ѹ��+�)�qXYz�p9�g���pH������E������{_������_�U+������r���sv,����ʍ��1�ශS��}�;����˪���㎮�����&:ȅ�GTn����s�(�|����R��FY.�r��/#�e����u�]��fq�J��T�����֘b����"=�rH���8����{�s��Ig�6���C<3{��7y�uP�R�ᙺ���驺&Gƨh"��{3|s��V9���J�n$y��ohmG2��Q&.���,��R���w^�^-��_����ӑ
�h��W�u_?����FE:I���ڑ�RoRȆ<���������:o")C2�im(]����u.�8X��>�>u��r��Yfoe��|&������������2�G�D'J�5I�tPFBF!���+���s��
���˨��B�F��N�mڕ=v۽|�A��;���K�-<0��u�B4R_4޲ɠ<��0߼����~|]��f��g�YeE�RF��[��=��Y�5䷺�ݻ��8����jCT�m��5�0##@�&�V�[��(`�LD�)t�R^ 
�(��ax��a�	��I�a Z~�җ��#��*�GZynj'��z��� �sSʡ�3-^Y�5y�@�T�-AAX�`���`����F#���'���"�&�:z��+�_=Ќ��>�4Aֱd�$>N�뼧ޗ_~yM;IY0�<۱��̴'�a~W'����I�-4�R�%S?�m�=��ځ}�;���,�Prю�<�����!��GGaO����e+�7;�;鶥n�b�n�IYl��1
I�44�Ҹ	,��  ��0���LRI��c��qۼ��ҡL�=�iJ�Zz�6�+ږ"s��ЙH}�K9����"S �3�y%�CK�;�2<�H���MG�^�A�Gz0��XSv ,��x�Q\�s����wuJ�/�@o��G�},<j������r^��P���<*$픓��͚�M>�eh���T��!�cr�vpx�+)�#�krj�z`rGڎ��#�јJ0�f��e���W���-����ѳd��<g�;	Yi�1��5��2�m��Mj�E7V����=Te�u��N� EG�n��^Z#ۯ�1�s�!�F�Y��+�mG�l)!e0���M��=c��ԛS��b��iR��~�6�+�� ��3�5�R+;n�ƀ�ι�7�SOr˅<���,pt$���#�6�Y�]uv��v�*Wz��"Se��J`��=w�9��� ;�F0$�@�y��<}@-p�\��c�1e}g"�VVe>u4�7�Mr-���:�N$�r�D��W.��$7m�Ά�)
���؛A1��0��Ns���Se�ډ�����p��@Y�	�z��IS�a�8�'/來OdS1��yc	
 ��bh��)
����s�7g�kM/D���تe�H ɟ��
����28�3�"vR�-M �1)�z9��:`���&�5u!a�#?� J��S	�y�Mʇ�%��2v����>�g~ӊ:��\�18������I Cd}�[xy�$<W�|�Z��D;��`*"�::[N�k���kȼ�N$,}O�4�}�EdA�.�L��MG&�iG���d#�#'�H�˿Y��Hj��6���I����)��z_~U}��<������eE1$�UQ�껣V����'�+�1��RbG,��u��Έ)�mA^��¼!J�Sn�ƀ�3�88���C ��+�O�NP���w�S�OR-��l��c��Q޼�>^����_9�%���f�����H������e|e�1`���2(�+uhc)�"n�A;��ND~����M��fY����Фfݝ6�����ɒ�4	���v�g?�ٕ�������-�OT���jowR�f	[DV�&����|I��@��\����/���{���H�I1�Sz�����lq�"�^��v
�Nj�l����D����ej@��$��֏9B�@p[P��L�Ƃ��k2jP�ͨ@�"�f��5���Sj'a=#g[ެ�va�F���(`�����w� _:ʦ�M�wϵyW��I��Y�,O.�B,]�3���a��ܽ,��pS�\��5���d��g؆NU�f�+W�2~�c�'z@����r�r%����/�W:-"!f�;鶣�j�^zY]��ƕ!f�(�$����(�'0��K�6w�e^m�tD��WRs�>;�g5���a-0Gm6����w�24I�d���l3��(C�9�4>��@�q�4q�F�$r�`D�I�	�	��&�a��y}��C����i�O�c�-�3?e�Z8ᵉv�^�y�(���	��~�l:/qcH~�(=�J�=��<t��j�������E�9^��\�$PgZ���L���S���������Kd��8�-sF8��IX�8���^_��:\e��`����,êG; OG�V31;s��A��B�f=�w}[�X�)�*̓y��R�T�NLq=C�d	2(�#���}ϥ����6�*=ʔ�̓�����vRƙi�43<�����h��l:�4B`��9�b�3N�A�ªo��2va�g�Nt^�]vY}ެ����v�au�<,��̽�y���oR2Uf/-ԲgZq�)�4���7��wo����o�SjȪ����R�-��ŗ\\A�HK�������Uo6�Q���B��,�]��K�1mg��{#�k��z}������[�vқ$G2]���el��?=��	6�x��\��I0�m�E�<Ü��.���څ���I:�\�����Ă&6=�V&�xk;ߺ������Q��uf&���x��_P��6{˙�l:���t(9�q����rH�K��f9��<�|�0��:gZ�4v�y�*
��� ��'V��7�[���=�R��"Lʶ)�tT��R;�.`��d�l买�3r��ޘ{s�oԼ�!�! *� X9 ���:[Jى�xq^���`�ƞ��2�6}��8U�tF�����y�e}��J�y;[�����{�ʪ����P�)���ző�N��7˪#�dg*�8�d���j_��K���2�7��׵Y�@��o���7��%g��Z�8ȧ�֮YQ�q�RN���˃�wY��>e,���7�_�=�s��I���_�ř������ʱ��\#�=ֽ�5�{�p����,�#^�7���^�Q���uݵ7����_s�z��J?;~d[��ysw(���}������7���������q��W�=�g�{^��o|U����~^����-H�>�T���뙈Rt�vE��Tzy��T�T\���On�f^��� ��i��Uy��";�
��f���\8 �l��Yv �}�Ҹ�<��@W-��W���@��
�u����6����&�
[.$�5A�Gj�EG���r�-	�q���:  ��٤��O���%IW��SY��a�w�xy.>V�2���H`O�i �A�-�6�Q�v�i��e��Y�p�+��LG�V�)�NB��\{H#uFxy�ic��MozӴ ��� ���߶A���_�����x|5��� �n ��VG���� �'� {Q�^Q�� � ���+Z(^�4��"�)���>���6��q��Q�S�g����	��=�	D¦bJ[�q'���^V�J|kj�o:�o��ָ�8Ӑ��0b����L���1J���X@B��ʞ�f�HZ)���Z��ҽduv���S<�Z8�]�ـ��  Ze�@��g���z)��S{hҖ �$y${�l��_G�kSI)�����ٹ��)��Ճe��v�yhO�#�b�}�#G1��zʫ�_;5ˌ3|��S�'c���T�dG��_�	d#�����6�7��A�>�6���_��}� ٻ�^�dC����ЃM ��щ�lDC/�#�ZG	����z]C�����F1r`��ɨ��/��r���,���ζ�:�U�4f�)nR�|�ì��A��C��!y�g��bȪ�<� "������=u@6�+���s193rʺ�{0�M�:8v2B�s�H�� jsC $�7���p��$}�v�瓞��͞.�D�k�:e����n~)�G�=�G}�sG��ۅ� K��=����̳I�=�:u
�y
�\���l���]s�����_Y.޳��؇F��ќ.�����U���m��e4bo_O�N5�2)@X��6ύ"�p�x�����4�BuR�b�Ƽ���K��+i�j^���B&�$ϖ�qf�3.ލ<�[�,�|�a�+;,t2�b_/@G�+�^?z~[J�Rۂt6D8)9�d
��9�Lk&����QaN�ќ�mK���t��l��0:�A�1�Q��s�Z���K=Sfٞ�S���:�2"3�m����a4E�s�3ْ��b�lY�=\�)�>��M�f�}{P�a% x[�1�~�I[�65me��Mu��2��r�#��(�rl�@�q:RPq�c[l��O��Tt�y �t)�tx!�yȩ�zm�z�^^Ӱ���:j��N��@}ԕWk���>3g(l���վ��x�V���ݵ��|��G�{�x�-�H��r��	�ȱ���a���sS��i /�\���V�t��3�gܮ����)WWq����n�5i��K͖�T�2�E�� ��H�[a2�l������n�|�y�hT����C-�ooGeݚ {�Q}�V���Vύ�m+���뻱�'��!�0{��G��MJ��f�y��H��V.�.�NCHE��L���sc��C���hz������U�b�:�y��[�y|<Coq7��� g/qHe=���֔]�u6�t���_�a&�OGǋS_u 4ʩm�#�cm�|�m�^lmR�M%q�Qy�>�Ur��Zu��ɮ7�M6����S/fKJYCO�ws��-J��I���t��@ݼu�è�M Ѱ���𼄣�^����;ŀ�3�(�}�	 �I�'�4�W@I�wI����|̓ZU�ɜQ��I�5�I�to���3�\�ZꦓQeq߽�C6��\�<��| W���g�^N�����H��>������3��3�2fz)�,7���B;��c��Ͳg:�G��VH����sm�����Y2P��#�u�	����n��YV�<���\�g�:o=��;i+S�6�.���>쥗^^^���Wo6��"C*%�O�"�7Y���B=���MEq�l���APdd!M:�x� �I�i���R�uܤvel���m���4<�[b~�u�ݣl{��KY�p�2o������ex�H=�{ϻ���%7���W����r�a�(�}ly�1*�=���O<��r�CO,:���!:�<�!Ǘ�NxXy��Qq�#��'=��	���G����GU��<�^er}`֔�U��gi�p��m�K2���Q\��׉�����u�(~v>���΃����G���Q]��(*e�n�3�kaS��9��zSIІ�RF�~W�ܿ�]�v�2�=��g�(<�H�9mp;O!�j��k�Ʀ6������9G��`%�¥��4�T6�+�4Ǫ�yh����p����<���=0��(*�l�=_q�թ�qd��+�Kx2��^z1�*�
@��m���?k� S휿�j�+�4v_|�J�FS�t܉ԍ�<W/�Ɔ�ʪ�$	C��.N�&i�sDt��I�!9��䷭��Tf�H=͝9�Av�4�R<ש;Λ��Q>�\δ6D�*F�LO}�3�.�ȇʿ���ʢ�v.�붔MXy
�R�i��T����f�?�EU�l��f��n��F��C���t),�X2�-=�vj7�T �x�6d��)]3?a�:˜�F"a,��r06eI��Qsn`��}���M^��\ٕ��毓M�������x���l���i�8�����;솰�BU����꥞���.�[�3�`���v��WC�ŵH&���!?2��Rީ�5�e���D(/o^�f�ɐn`�)gᓷ5���Q7L8
kG��hW�<'z�V�1��Va���*t�^o�5��z����Zz�ǻն`��!c�C�`��B`�v��w�4��8\ډ�O��vԗ���5�R��T���k�^��'36�j�Xz/�ͷ��yw^ `l�f�IYȅ���XT2�mQ�J;`�����.���Us�W�s�Q���=��K<�<�˾7)��`X��-�T���yS���XYm�R�m���N�����q�{\���
��7�_NS�ԕ�R�}fÝ�4�S�6��@U�@�pu��xhd;�}[�l{�P�����������H��&M)\��;�;�\�n#�|M^t�ގA�Wf���È�@H��d@�(�#o�<*�˞W������i�v�5gF(���������H׼��%�H���ԉR����)��z�|�xf})&�C�&#�2,��3ux���~ą,z{Z_.K�%��"1�x#��׆x::��*���-�j;����g�ч�|�L`������-{�t����������^�^v����i��fC�lcX���5ӱ=Py��mC� T�M��<�{@�����D���:��rӲ[���	�*�:��ۘr��b��$w��h�N�����K́U�H�R�Q(��X� 8$32�Z�ܔ����ډ���Γ��<D3=%Eǀ,?{8J�Hj��yrK[el����_��8��9f��*�L�6�	�|�̿����<q�L�Ԭ_�-�u��ӑ�y;�Ǉ���L��_2 ����y����"�0��g�= ���d�2$)/fG$ކXؔ{2�i��ց�Ѝ��Y���t~F0��F0�sᲝQʲo�D���Z-u���)�C�z�q�f"nsX��]���N��J5�\�=]�N����vO�񃏸��e��}��o˛�0����>c
�"f��y����ے�ZS!�4r��1��K��;z��Ծ���;���N�ep�l���06 �2N��s�ޙ�x��1��ڐtC�F���s�1]=fK d:��<�lݧ<wN�3P��7��{��9���Y��[����`S,��rJ}c��*~k;�� �E�<�@LK��ogs�9]���h�p�ݚ�ŬY]��b��S��b4���
3�yK�/q%���p̑����قa;R�������C�����s��)����M�(�E���\#}��x���+�f.�\Q��{]��K�qv��o�٤mk�V1V�����0M��E��ʁ_G�oҶ�A�@�J��@Z�4�9Z���G9Q�q6Ԍè( u�/:8w�'�N �<�c��8��M8 �."aq��<3��l���|։� �N�y�>�Kg&n�m�,��`��g1�\�O5�/�Z9wm*�� ��[x�#��޲�=�2u��)�M��-/׼��f���I�wR���z��,���a1�u7ϻ��g6��w-�,�ћ�c��+d���ZyV��BpǞV!�xk|%YB�\G�I���7����^c"˰6CM��PvM31�o�g�at|����:�<Z�"|�9��Zt�l#�D'��[$�o8vGy�����jm��V�Z��r�J�{<ΥԢn�G'�MV��q.����F�BՂE/��Y�je����%���	�Z4���l�HR
�;��d��b�x�ԋ���
e�i
��ሚ��u'nR�����*��!	�L��,�#O�Ǫ�:	���.f���!�����(��"y�0Y�����Vy�gJ�ν�v} L/ q�@ZA*�j��c���ӛ�3�Nl��
��S�M����I~<T����j�)�ds݀3��9c��@^0�����<�z�vo���#kۺ���/�x���Q��G�͔!��Q4I~�Ý�hrΛN��&o��48@���./}=�FK�W$��2`�]����5ǈ�D�n���Qb�����(��i�Y*�_��wae(:���10�1:;y����%�7t���6�^	g�Xdo9*#Q�H6�'Jo ���e�3|�������ID�w����*��|A#V^[�֬i�=E>c=e�G�d4#�HO�d��+���H\�F�3�?Y��I�,���r��W�qi�7�� ���I�T}����O���~��
��4���D�4:��‒/6�#
�y��W!O��Y�L�yO�"����]K�
&wUV�sN(W���,MFZ� �I_����nϢ�w��.�Y�h��(s�� �������<f��krR�B���Ir��]f�!�'uj�-E��C]���6�D�d��y�3�0�e�^H�	�i�k.�"=��R���������5�W�ꍆ�G#2�q�@#�(�
�����O>����IyV����/�sv,�]zCY�Į�=��5�l���v,C];���k�ޫ��ݿ�X�S�۷,]9�w�]�z�)#��V�ާ�u���O����x�.�k �' =<y���(ښpX���F��0�����+:��l��9��q�/G��{zB^�e0 ��y��ڨߐ�ᤍ��5q�|�h�*Cc��p�+�_YS�)�����G���_[����r��W�w��-u�e&�vl-�ɦ$ o���똆ּ�it�-�Yy����6 �K@�8=s^#X�Tg���uNF�u���x�V���ٲyg��vv�j!��H=�G9s�F�q֗��מg���1tm�x6�=f�=���>ڈ�Uh��h@�cE�\�Es>5��d�6��׸�d�)�&o-�}��7]}]Y}��F�b� 7��I^w�#��ܴ�ɚTO7�:��5ulUd�ێ������+k��)�]U���`ٽ��#��1�>�����7����l�t-8���� ��.Cs�-�sX��<��9���9���9���J��s���΋���7p�wNp�k���X��vG�S�g&<aeW��cފk]+�p�/K#���;��v.KW�� 힅�H�[��-Q�2@;g���� �������}H)sO(e��j^�+�t�S��T�S~�`C�9����m���hc�F�����!��s�񓓚���P���t�t\��Ox�?F�R'R.a쪰�	�
�>�9��P��r��BR�/��W9�g��L��z+p��ٵ8����l$�E�M$�ҟEu�X���ɯ��3�`N���ڵ���f��cӞ������W��51���+L�.��ȋ�&�W�YS���6�M'{j�����gG�������ѵُ��FG��ϋ����22��rѹ�+�Ʈ*s#}S���ҳ <����#ӎ����Ԁ������p\嵾kʨZ8��Zߞm镩�:?��=�-c�=���o����^P��|x9�����_s�����◔O�����[���/�S��i壧��RM�T�E�ݕ��}1�����+.*�����A<��Y�U���Ob��[9�����5��.8���=�G޻\�����u9��Ϩ�r�e�+�����W�Dy��Kʼ�C7����s~e>�p�受\Q.��r�IO-���?�`O.��S~���+�2��{��i-�r����*QF8i���ASB�<G	ɝ(Ӥ�@�Gix眢��WIi��	����(m�Rp��^��"���z%�R^F.-?��K[��Fc ZӸ5I;�)yfy����:ne��i6뙤.>�hQH��Z)	y�;ë��s�I��ۿ~�n/��?M�5/o��^^{wM�4��o�`� l�=���f�ⓓ�w����Y[�ۛn�������?A6e������`Yd�[�]]�MZ8-]����������f���u�~`{�Ǻ�ڨ�ꨃ��5p&���g+��������c��j����*W_uc�zwYz�`��vޥr�����yLY3�s���_ d_ ��ṟ�ԩ�g�~곧G�J:W��O� >��{����s����i�X�K9��������r��.w��=ˊ����W���RC�r��?T~��ˉ���^yU����˯+������ʹ���< ʲ����%���\��?����p×����e��٩��GE}w�2D����l�zh}��k"\ٳÃ��y�3�<��K���R��&��c�\"0��~�`�����Hx�AѥaC����%m��Q�(��c�X�)`Ш7���8R6���Q<i[T�*�U5%!<�^����*������V��G����V&�Y�M��x	���X�`���)'����=�V��P;�n�Z��md����&�j�&i;W�uۓd��G�M�ݜs��kV�6�����}YY�g�tbӚi��y�由ѵex��墟~���������5����\�,�?�r���*L�h�vuY���|��g��ͺ�5\0��-k�z��51�p�bZ��_�l������-w?�e�}O�!�.e(�z`��� �O��� �O��g?� �綒u7�ѵ���^T�������]���!�����]C��e���e�_Y��'���M�|�,Ͼ���5�]�>h�p�w-k���N	|���(�_riY�bu9��U�r㥗��Yzw�;�����7�0�X�멋�n��M�r�Me�����I|�?���?C:�|�!�Vp������s��h3���x�� ��FlR��|�$O�W�!��w�[l��������Ȕ��0��>�N���/�eqO����@a���d -FЊ#��O �B�:���@��$��[�v3Xu�޳���y/_����)�*/~�+��4�Zm��g[�7��U��� `0���هt����n޼7ս	��C���RF��π�1,��~�r��_-�̍�����pV��[��=�-RS��:Қ&h�L�9v�����7^�����?����}OY@���E;�G�3��7:����.�|�Y��|�K唿zz�L�'��2�\��q��3/�tۉ��NЍ.��q�2�u���˴\�SA2�+�jkG� ��E�*�8�[V�,���6>үr����o��51:jr�>�i�U9��/�^�V�@�*jϡ�0!�)��sFσ2�I��iD�
x�.ɫ��I�$i	/�}�@R��dx,^��k����}����߫@����U�2��;�!����wʷ��nYe��g-I�~	V���y���2$*�����I�b�������ʴ��~�]y���@Z/�e���%�R^���o%����~�Hڒ�V@�n���6�� �E�ZCAˣ����m��~I��b/��#�:]0������>����T�!o� Kv�h%Avμ�!� ���e~�ueAO�^���HW�*Oz�_��.��U�M�GҬ5�@�h_�j�x���~gy�#O��ۓ��Ը-X��t�)k~��)s��+���E��O�~@��vd?��H3��i�l4 [_�g�.�ţq�����T� �8����jW�zܔ���B��{�D���n�W�������b�d�(AV	'�~�ԛ4�|�)a����q��wݭ<�Q������}Ua�i�:� �����:g�ّq9�{c�c���<QCu��t]���=��o�Nh���21M	]��ǐ=:����,��k�,�|�0ԓ��N:�<��������>��\^ӯe폴|�5T�w-G���O���"?/0��XV����N�o�.Y��zc����¬^���������?W�Wܑ��-4�.v�qa9��ʃxT���r҉)���G��vR-���'��qbQ"�
�����	�8��66b����ꄧ�� ��{�e[����q;%v$7I=��u$'�!��N��� p��X{����(�z�,k��]&vد,��|���=o��=?�qKq����y;�Ѿ�1�5���\�l�,�_VM,.�{��y{E�h���1B��`��2�g�n��D{Nx���Yd��g����z�-�gS�#�p��[�7�>_�P.��e�S�|�Q㰘(?9�Kg]ޑY��r���x��*9����d���4�g4z}�h(�x���jd�����Ct�ǫ ��}�Wjh���z.^���\�)����~FG��'Gϥ��%(i��!td�#�z����|���,�}��?�������<�٧����;�;)���]S��J'�Ri�W�@�lc9�uĈl��xA��@�`��t���u�}�G?�����7����{���r�{a(hԿm�%�!cmiD�����9�\{��oS>to���A�`Ɇ,�������g�Y��ݳ��3����o�[�r�9��?���-�*_~mY���l�4����� ���eh��,�y��k9�̳��)g�uv�Z�����|�̳�ySuo|�����A�?on8��)���K�Z��#�n��$���ϒ�6f��ЭM���1�V�Gq.JFk��nh]G8h��HY�r�zXz�h�ʇzh�2�,���e���-B����90b(��rP�E�7p�"��؊c������7����lρ��{��B@Z9�^?������i�DYvˍ喛�+7.��\s�³�c���K��7:�2�'�T.�Ɵ�#eW'�gʱ�,-���cZ�by���D=1,[�jY���˂�8������rˍ�DYGBh�5sz�'���dAޮ�H���.=h'�l��6iC�#}��z	hy���\�d�ϴ��$���-/����-nثƾ#�J6��8�G�麲i��o}����~�ߔ�����e��L4i��8[o�>���8M��n���|[RbL����]y+���Q�z��o2�_�S�I�5�J(��	=o8BBe��W<$. t�ʟ�uJ�0�fX��X��2�45���<�����Zn��ZG�e�]w,_=�K�kg|�|�k_*_��'�W����Oʚ�e F㣭�SQ���,+��7��Iga�\u��S9P��*�ɮ�N振~�|�+Q��~.<��E=?�ʍf,¬[���mO�����6��:Ѻ�*��&���FFG�W�۩���Q�#r����bKd���2�gv��:�����<@��$ZSy[Q�Y�-�W�.W_~U9������=uت�E@�\�2�Ɛ��'�(.��I�S������ N�-�:�|�ed�6�_��$�c�e^� R(d�-}e���?9��|�����g�_=�+��\���rR�:e�
���F�Ԝ�Y�!u����1�E%�U$µ��?�O�39uE��8j�:�Mᐽp�QG���b�@t����ᛴ�G[�^@6�- ؜�S#̔_ڧpi_wDF�)3��
s�S�'{Ɨ�Z�������u���z�Uc;[e(|*�����)�Uqo�5A�V.���މ�l}���r�
���G<�1�k�ǐhZ��i��O?�O����K�x�u]�0��#ep�`9����o������<�츠�<���������-�֎�7��#�̳�*g����o/}UY�h�(G �D���<�r��M����Kdפ�l��k[�՝!�g�(�"�\Y>��O�k����3?�q�k��-���i��|9�'���e��O.C^��\]�	��v�i �9�Po�!�A@�^_��#/>4n�����D�x@G�^�my!���O��Ou'�7��@���zl�ҶDCS�r{�.h�e;�v���tC����?����?R��9�wv(	��$�j^t�����N{�w���e6��m���hz�!���g:j�!��"vM�ML<��Y�r�ˮ�U��6v��`��	 4�_��2أ��
@h��n|uIOD��_�4(	a���=�	�HlP�!p��`,R&H�#ce`�Ϗ�B�.�t@�����=���p��Z��)+�&�[�����o}��u��_���p���ܬ��/�>�� k�os�� ��A����� �N�=�� {Rخ Z���5�|��-G=��I�}�6�V�s�B�d}ܗ��XݱN֏ҩ&�z�˯1 i��d���]��^���՗P��nl�M�7U֨���Ǟ�	��f��H�MT#��#qn+j��f�Y�,����pC݆w����d���3�������ٛ�`���pl��%y��{�s�[+���*�X0�~�����+@�/ f<{�(�tO��������Ã_J$�}���<�6I�'�vhU98@�;g�Q7	�|�}�x�'����e����կ�px�_+?��/��_���`�!�^���A��Ų�NYZF�	dy��H&�'L*���K�;�\{�%!�w�?���
����n�@��O|�����d_ �� و�UG���09����� ��� h$B7t�@�B�7�,�� �l_k�D�^`�)H�����[zA*��O�������@�o}�r߀�LG�z}S�̒����U�6��"�f7u,ɽԵ<��%A���t�?����=���w,��Ҷ*s�#^^��G?�1ext�z�c�e���]�����D����Fu��
��䗼d	��L5؝�\x�0�p�&b`��<X`�Q�:3R��^�l�d8:<<�����
��{7/[Y_�X�0/�#>e�̭9��V#6yӉ\�=j�&R�q�O��JZ�h�N�!� �5���v<ᒚCP�{ scyc)맍�c֖:ez�����D��}/��SN)o�ۧ� 2��*�
��y��9�yN���q�8�M+�l�e��Te�:�(j��)�$en���Ee��yUv�i�z����g����E;{f��>|¶g��l&�a��C��|�z��:R䅻o�����e�b�.;�V��c���Zl��c㉎�� �ډ�`U�0���49��x���U>�r�}�)O{���p-��/~�u�o� H��}�|,9{�Ɓ���5Wە�*c3l�9a��G�͹i�/f�t��(+F��iBxK����^(蜨�� � ��%�7���Ԧhf�������thy�}���m��X����2:f�o^�i�=�y�8�M�JQ�[y�-���Q;e�]��O�2�&k뜟�<��\<Dg�t�
��K'qZ���m����'�')g����<�n�&��9&m���@ݾo.v����{�=�ڽ~W���'�T���>����2MP�(�hs��xe�b��8�Ij?'nn�\�\Z~^�"� �kQ&�#OF���\3��uHP9���=�y�r̃N,�;��r�Wt�����_�����z#�2�h�k�'�HٷS�����
�;�G9��?��r�1'���=��ɑǖ�9>`^{�@�Cc�J���l{`���~�Y�Β^]z�u�K���ܗ��g����lv�tʶ&�U�K��J;�<u%��\j�fϳ%A�Ftg&�-���dg�m�Qr�3�N7���x��2o
o"u�Ǡ3���`kx�����~?�Py����LΩq�-( Fʭ'B��i`���e,ҳKA:�!��e`��8
#���l�L/`���jy�ɞy�7ˣ�������>��^��E]������<��V>��/����gQ�W�!M�2��vܰd�ɖ#e��d���ʺ��Ǯ>�U���/}������|�_+�}��ʂ�$��%��#�ز�](/<���ǟ
��"7��� |KS��:��:�]��۬�c��&z+ɝ�e�֟�W�N-ڡ���W�W��G^UGy��iO{Z�Ї>T^���]w��֔�DI��[y�Ԫ�:��D�m���{Q{�۩]>��ِ) ;�.j�6�T��V{u���7-��p`�����oO��:\a�������R�P��_���GO+�x�;�P�J�PAm��)H��p�͕�$a�Bq.-�n��D���ty.@YX�&'9-nQW.t`9+@�1�zDY�x~�{�=#\k>Y�ܲ�|�����J�q�lt�t�<��]�y_���?d�[��+��������׮)_�����Uy�[�P���O�������o~�[�ǝTN}�K��ǟX��	��Z��5H=R'��0��NOg���i�u��( �M�<���gM}�Y�fj���W����r:*�|R?̣#��_��Խ�U�u��I+����aj7�;A�E�r�ɱW��t��i^\27c��NX�4�hW��xf��M7�X����w�� b��	���"õW��US�
�к
vV���v�](p�7x��������Q��P��Y�&�j|�A��~�<��o/� �i}��/=HcN���@_���3��
��d��:�/�u �կ~�\r���>��e����͛gN+0B���'��S}I9.@VZ��"��>��H噣�߹r��0	�⭫���|Lx��z
����=O�q���QB�w�����-Ѣ����z�-b����^���ڡ�u$�����j}����h�<Yߕ���l��˯��~�E��0���*�1T�;w����W2�q��<��/!���L
}��[������O��� ������|��D$�K::���Q����n+�,,�}�u�x��C�ʀ�څ��U7�ޖ��nA#I;�=S����c��y�9Չ��ΥAF:d��3��ͅ3�2Ta���;i�{�dm���)�u�{�N���i?/� _�6��F&��g'���=�=P�bs��ٸ�DQ�ݖPJi��t�g�&�Ɇ�ʦ���;�k�g+W���`�;T�޼, ̜�-Dk��U����˷���B���yk���f��N�GA)�*����p\����Rn\rs�MS[��?;�Nr�R�,�����'ۗG��^t��K�\�Q֙8I������|��t�%��	�[Zw�:"gL��m�(T [SBw=��r���+GsL���~l����h���s{�:]����gZ�4`Ai4M�4L������a�RQz2!��:$@����v*���:������򶷾������@�Q�U���zj}���x=���i��lk��{�S�u�\��i�X��m����p����e�ؿ��}��2��w%���0͗����sϖ�Ƴ�Y�G��%˹��2:alkWO����7�<�C�NrI��iik^}M��ƵZ�9yL�d3Q更��o+�.�&�	�5v�c�t�\+��C	�YqӔ���駟^>��V�ao^��[h�^��d�A�8NG�Y�u$|2"���^����!�kƘý�|�L�*G��7�W�鑏xD͋���@��5�����e����@��I���c��%����d�1[�.&#G �|~rǶ6�Lʿ�2v^��ϛ���O��	��v�iu�H]�`ݭ��[�RF�W���֎d�^�d���S��ΔiNG�w&#˅�v��:��<h�\nM�9�	���\,fچ��}��޷t�o<�O@�C�	��o����Yu�׻݂솨�r� �p@y�����cd����2P�7��o:�Qz 'A�=�㎋k���' ��U�v�u��6����7�/&�V��Z��)��i�595�>��4�=�E�T9�Gz���;S�Gґ���H}Wع����� _m����7$�u�=w�;Av�������vv�|�����^ex��3:��X��,���.y]��_�o��n��QE�Y��� ���09���\��������o<m*1x�����{ʗG i�G��dGen�_�1�i�@�Heh�ܳa����ׄ�#��]�d���n�����~��^�[���ɐ\�B�s�M9��)�lc흴}}@l
э�ɟ��8���6���Vi�O�=������cD驴��<+��P�L��0��F�J�DYF�l	�8Oj�7�� q�{�'(n.g�y>[jO��^�ކHǘ$ܔ���}���:�m	dI��I�Gl���y�ȴZ'�E���	,��y{���dg�46*#$켏����D�`E	V�x�BYG���&�;��f���t2rokP3�M�fٚ��:d�S��6v���e����+�el����훌u���G]�`�u�^_F�[�D�֚���1 X�C��m2�^zp�1�aA/��F������~��n.e��@�L�ӽ&��)~����t�B3=��R�M��&ۘ�r�'w��M�B{�u�Y�cQ:Y`
h��__�)�6�m��G����Y��Vi�@6+9��gj*�������O��]N! ���mOS���ϔ+YG����0��7�����Y���f}6��6־9��N@�B��f^
�kv������,�&��������<Sol�Ƚ�C��k�^|2E |��u�]0-=i�ٹ�PW(���m��(R6�6@e��W���Ӽ��i|��R�ie�M�to:���q6&��Җ��26�?u��Kk��aaO�fw��y�V�7��5�h��I^���M,������AѾ���'��rJ9餓�S��!�\WߙN'k̯G�~�u�λ�����EA6	�28CƜ����\�ۇ� �9J�ˠ' ֔�cN�J`@3���$7����N��4zl���:7�W�J���پi �@?lӴ��/Y�!�Y���Lr��h��µy�{[��D'�#hG��#	i����Srk�'�?ۘ�ٜ���}��ɓ;(i[�4��i!:���巬���N?�P��N����m$w�֥�5�4
J�(6���ɓ;(L ��o�ʛ��\�l�:姯��l [��0�!�� �������) �-���w҆)q�z��Gk!�����{��ɾ�E/�?3:9�'����NE�c���Imm���';mH>�[�;�'`ͽ�*j.p�t�/�4�΍%�,�`��L,_��Ε�rc�Lt'�ޱ�N��<����ͣ͗ϺR�v�� ;����J�W�\�d�o�d'Of��dt'��L[dQ�Q�dK����s�$�A    IEND�B`�PK   �N�XWC��)�  � /   images/093f54e3-331f-4155-80d0-fca9fbcaa25c.png��	8���?>ҡ�)�T�9�TBC�,5��A�(Kd��/�q��2r�fP1ɞ�0�Q�
���=�k�}��~�z���������{����y��{�_���ǣkښ<?���\�����.��~r��>9��"�؉���]���u���K7�0ؑw�v7����0�='k��-�;0��v��h�[�wN;��ď�?��
����O�h�O� ݯ{~bz9a�.n���(��@�n�OoF�������_��v,ȋp�qW,��!��U�Է��N_�W��+��ޫ�}���.}�s�����}2lTSr��i�� C�s���sJJ��i%������鮋��?�������� T�źȜǾ�'w��A�t�+��OhEz8Ϥ�/e�>���e�%���%O��'�3W�L�����TV^&�o^����{��b0���.+Ű	�~�8�O�m���z�K��n��矌�t��d�D��`���JJJ�a��8�]\o7��N���;�Y��Kxrt�
Q����G��jm$M�KBS�='{�VVX+���i6=�˯�hT��_�1g���a��p�ݥ���6zC�*��4?,V����U�\p�{�3xc�w
C���\�"��	Z6�{��O$�O�(����Wj%�X����K���}�u�=���'�5�^%U_��~��!a�@G����1���̦a�w��W���4�8�$,䄞/���v�G�����^�-^CY�	�S�	�n���!T�17�!~,){$'L#Y'I�c�*1��9H	���|$��~��P�M�P�?%ͬLZ����{�OY�'L�oUۿH�H��������e%���OƯ���CkBW���Ou����Ƥ�n=`���C�\������Ŕ����ORŖ� ���۟��(����򣂒WP0;��e�*m>���G]�
�i�jl喨4eX���[\Hk��������6��ņ�\�B�m;�=��U�C�89ݻW���sv�~7%�f�J������n�2�oQ����u���^ۗ��% �5��£9�Z��;��� �1����p�`�g��7�Zt��nf��J/���DvE�.�5�b�`=ۥ��"֛�����K��ͫ��C��zCq'�sN�z�N�����j&ӟ�Fs�/��!�;�p�ԓ��8�L�aOǆ�{�����BT�}��dPTbߘ{1�K� ]���`��8�6JqSV�K�O���0�`u'��oB-¼�E��a��+��G���s�.��/�2��|cB��6]�`�2{��TW��wAR>ڦ�ªIϕ�s��}�z+/��Ra@�;�b�.NӍ�;n�`y�O�X���V-M����������D8`y��<�D�Z�5����`ҵ[���X8>�Q�+�Y�m�L�Cp5~"�i!����a�
���	�MO�����B�"��2�T7����\A�I�o�}8�àq�`_�K��w�.N��<�_��r+���>�m�0!��	�?���c]dkjd�9�f};OA���HGX��[[�klHR���B�I��N�-%=]�$X�v"ɑ4n�<���v�{Ы����1�����m��(�_?�'t_'s��n7�Z$qR-g�}�����
�3�U�	�ۉ�Bk��c�4Ƕa��?��d'L�_�� L'@\���P�>���u�y�f�O��1;arQ�	$|I�KՎ��^nKɳ�4X�,D�|��"93��"���$�7Y��y�������@�N�K�d�ct���}u-�D��g�w35_��e� �2ty���dM��E�Uಷ�'�;6>���X/�I��>�ѱ�*&��7_�~7$c[F�O-n"Y�'������N������-��C�*6g�uv�����'z
	��r�/@B����p�\j>l{� X��P���z8�&7/o_qq1��w�7~Gg� �5��O�|��Ijs$����md��41��=�Y���E"��ll�]��wӵ��x�aΗ�����b���w�{q��lO��5ޣL��3ZVZ*���L��6C2�\0��`�}�^,��J�t��B)��x�K��x������$zU׏׌<`ۋ��s�.���]�J��ˁ���#�9�!@'��q6���$�����/%e ��EM���ˤ�(r�1��zI"���� zZ�	�����߾=JM�>����WW�e��Y���9m[9L�(�������[��K���G---����f9�1{RYQ��&c�.E}9�]�Q���{K�r0?��%2�%�:^3�YO����?��dH�UND�k�@ �lz����S�9��Fp4�����h�]�|/�5�_DJT��'A�����^AW�H������ b^��z�����z��efeU��Z�D"��e�wI�o���Һ����%!��k�K��n�^������rs;k����W�+���Ȉʷ��o���MI���Z�]��󘻕���w�C������FF�@s�F�j��[�,�HZO+�qm�n���@_�w�{����f���w�_��6r^�@�I>pC*�ӱ���q;۞=�)�@e�A1�E#I���+k^.uK���'jM?f9� 8�� S�@�T��.��w�=��U]dnI�p���{��%���kS_���S'(,�Q	f��.�����f�kn|���Q�+#��
 ����g�T/�����Y�y:a�x�[�%���*����f�4UQ@!/�2��p����W'Xk����u��ӧ��e���[��S��7��c}:[w��1��rv6�b𾿫�a�g O^k8��<���f�\^c\�s0���Uv��w�
ܲp��V^w�� ��;��?ݨ���MC� �M:�M� C��},\K��RZ�B�&� xVZPp���X�{��E͎�Ύ���S~�=�y�tWj@�XV ���<G ���ؓ1�;Zv���5���Ά�V��l��&Z�	Jh�^��kd����o������������{珰���6�)���i�,w�&o�@�X$Pڡ�� �4���Fe�)<�8��O�!*7141	u/6U\�� +܉i.��0��O� ƺ�:w���f?^7�^,sp�f��t��lhf������8U /���@����l�T�	�5��it$�ޘ��%�O)>������Y{�h���t�����	�m�ja)P<͇]����(wY�o-yꔧ�Z���x�[�'���<��G(�mm��	��X�����Rp�[`)}�ROG�H��F�E�8�3�	]��}��m�L�Z��k}�ES]�w�hA�r�����C��ќ����.�&��-uC����|7˴{a֨��fvXq����Ps���<{�#S�Z@�S�d2����U�%V��ә������q��������^}Avֻ�s��j��A� ���f��U�(V_�N��j���3E:�SO(7�|0��5w���P\ؿ.,<�<g���� ��Fe)�X+H$���4����F_YLb2���D1�_ל��.
u�ԩH���gv/V�O*����w���AS'��EA����K�W�"i�Ts��_Zzz �XPP�'f�V�u���7��:EvQ��~��}]i�Z���{��oG�+��C�3�p��HF?v����;<=�Ez�����&[���j�����$]�A~~<N���ie."��Je���]m�=ɧ<���B��p[��k(���Z�g�_ou��Cj��Z�7�]��:�/EEhV�Y-6��L �W�u_�X��M���y��J��z�k��/-d�!B��������ۤ�3�6hBU��]��4�,��� ��%���^�B	���������6�F���ă{��lp�őhF��Øq��~�,�G	�k9-WvĢ��p�@SμL]��.�bU�T�99b���}8�u�HrDq����\��j*bcku�M#�� V��Rh ��qprR�z�"��ž�AQ��ĵj8�}}�EW�#���}l�<&�8�Q���xr�wR��`��Mӫ�
�A�M��(ƭ���M���o�������)+۞$�ƶ��J�%%E�]}SR�;j���oԦQx�])== &8�����)�J���u�rY�o	���Wy{��_�r ��Y��=�6�WC��U��<�f�i"% �k��3r�"�zC�����gC!�,�J��b�~�����������n�	�6tBHB}��z�����d;����8GRdg�w�c@��
��l�����0YeNl{JJJtqեӭ��d����(�ȧ�����tl�3�l��vd�gS��J��I3����?ͱ���6m�c
^S��IV=T���ODy��t_s�V
	�]���+�}!h͟;Iv�f�B]Gը} i���4">�)tf����<4��:��J�'e��-�([.��z��.r�)��M�o �0d����wHGܚ�/f��?�T������K���k�=�����o ���>D������C�5a�]���+y��_�������9�f��*�;ǃqX�U�^MO�p��L_�6�p��͆7S��> H���j�8}�N� �V�5���ւZ'��QH�������9����Lv{�M5���;�]:m��{X�yx6�
�U���ꦭD�X��l �@�T�D�)�]��<*la�PWo���ux�j��rF��!�Ne^p����O�̸�t����_�YC	R4���&���JJx�Y�.E�ɣ��S���p�j�T4�J���қ����g��.�Q�'���E�'�Ν;WF�삭Q�f�j���1�6���ک�<�éQ� �e$��ݟ	Z�Ys3��@%�-bz:T�)^�/��~q��SfK%�/��^6�ʯ�$�DY��� �O�5쳳�SF^Wm�+$Q��\n�$ �k��#؞������,��I�#����@+p�J�Ȭ�>����"̎'�~�����o�ċ����GX;]�z�@�~���&_֟˝F�49��Tzϒ�V�����Y��s�3�g��`,�H���k��yl�=���9>�745M����j��Ry��w�TB�M��	~�[� ;��`�h<Zg��~�v/wu�4����6Sz���J�$�ZҕђH]�t	�訥#P�>]�?K�����V�Q�;-���RampX�Ř_ާ<Q�hߤr���R��t�lΣ��D�Pܪ�=劲�|�������e�]��cl��֯�R`�,}�6]���.��Wf��\+x�+��W���s�Sk��q,���Xwi�Fc���}Y���l(��+��O$.i2P9ި��҉0r���#�h���ȁ��co�M�͡O�0)�J�[��� �������𝮟���S0x��1�a�tB9Ɛ�`�G B�KT��Z�� ����d�|I�u��]jDؿ���*@���v;�i�U�2<T�}�rjk�e��i��������Q�+Aw�&�e��=|2;�����R\Z]�:�$��@�%�1�z۸YV�(P����Ŋ��],�|M�G"*��q�j��r�J��,y�k��䐐?�#������������&Y�]^U���3�8^DO,y�w��\����>V�<߱���(�@�ƠQI�k�,�س,//����,?%��1��˫h�g����Է�S�Q:b���n�s�{�wͼ\h|�"���I��)�i��+D츷��� w�Ә�i���kÈu��u`�����$���v���-T��T,��UE�K�X�Q���g�P�A�fؙw��a2@_��5��8�'�fyՅ� �"����ay]>�H��'���$��[��
&�Z��}��*!Hu!�s�x�h(��ݾ��. h�P�s�*?��_�u��Nm�ݝ�~�C�V����������W5S���7�x�L��h��TE�|�A�����A�#���'��ݓ4[6�Uno�vB09;���L����;��q����d�I�H^�77��7o�G�z����O~Lf]g��&+�k%}pM|$��KM�'c�Ck��Z)G��B��Nii�E��ih~X��|�~v�l�r�M�����J�p�sM����bta��I*���f�����\W��,�c+$M���g���Lk���6;Zq��ɓ�c��m'&&X��o��[�VL.��dc�)-���%���w<���n:���R��l��H�cW��)�M=5��KA8�{��Lj��r���s���$�}a�֜_�  �S�O��w��>�ɂ��B��������5R�Ua0B��[�2���Qq�9�#�o߾eZBlL��o����/ �����������X����gO�?�7���_6����j����H	�xr�M¹�-g����3�ƿ1(ZӨ��i�#�X��IYQi��(�@+h�X~����pG��E��֚�(TU[�ԂH�}���S�F^��<?k�PEU"=[+~�C#,�\����RqQ�M�\�O�0�
){Z�5_������֞���V�i��mvv��	��bd^��I�ø{n�x�|��333:P�����A�p����x(ӎ�����AqmN;UO��	j?p���|`�g����� 5aW����'?p��%o�
MB��ϣ}�`FisؾȚ�7����nM�brA�
�	���/t�2¼}��Y�0a}$cIS�o��t��R�A�(�6���:��� �<J;�d�X�bB�xZ�ܜ�_�OhP���=�oI$-�p1���-��'� �"�(�U�	]����^��9hbs����ؐԶb��:%�ؖ܅?���A�TS"�n�i�'
�P76+=�-GRr��fjs�U$�~0�&��X ��KӻZ�>h �q@�=������J�λ:�A	����
b�<� ���ݹ�_[|�E�jf�)I>��� ���U�h	$?qq������\$�[�W�3!�d�&<f����Ļ!������~qm ��6|���TLX)���<��Ьw�?�-�x� �1 ��!_���C�p�r�~�M})�y8�7� ���;;;i7����h���(TPAHK?��꿇+�U:�|R�(��
>8?]'˞Kwu�12�~��Bo�m�C�O`i�;��@��:نJ�V���#1�!����>��2wfD��t���^��s���0"�Wh���[�m��W���-��!�`��gc����ŝB! ��84s�*��IQ��@��8Ȝ�995iz�� ج��\ޒ1��o``u���o�><���[�hȽ�����M�v�@Un+|��Ǟe��� l5�ѱ1���k���aY��T78VFy�����/n��R"�k߹s�#Z4�4�R���c[^t�BF�wS|�#I�n��Ѻ�)
u���T'S�6����w�0� �����/��h�>nAd������?mP�}���M���㝅�@F��&���{{���e	���Yb�����A96�	��='kYq߶נ�2��7��(|]�_��J5	�Om�����r�;G�����fF�6�]��+֘��}�H`����у������O��(t�?���̗���vh�
��2��/��
Ƚ���p�߫�NG਴CU ���{"��`������z��7\&;{(�t�u��V���D��+�n��SRI��R����n��}��V�翐�����2gA���r_:p��(� h���A�@�5T��.�4Y�St_��k�ׯ�����`	���F�s=S�a@_���ͧl�����9�k�f
�{2��Z)pڄ�"�<�ޅ>����% A�
��i�t��rmSu���QI8c0TT���w�}g�w�燼*�
��]MG�A�(�q�F��IԂv�<'��y�%l5���l���b�V_�P'�K&��!r�^��%�}�i�}�=%2���Ջ]{_dgqx�>/���TF��=���+��z��h�s�n���w
��B���u�:dt�P��x:����ms9�k!�t��Y��n���c�p��ۭ���T�is�-���R���w�@mԶ=�_V\�x#�[�-����������`�ݸg����@�b˵- a���}1v�bon[�]��_���&, �b�a�7�I �Љ��	� ����
����䓟�1j A7Q�Y���F���Q�(рN����goG//L�a��� �,�g���:8�uX��7����{9x[�?<�z�>�/~�s<�?��m���Y]�5�/L��<�ǲ��o��oT���u��������޶G�8K�6�.�f�l�W���t��Z�~���~�F�����ȝj!�FQVgdo�S�(��(���y����e�D}z�CдI��Kg�˶�I��k���/�������ہ���@���o��ÓǠ�`y���
����}y-nVm[qLbM�����A&)�9����I�������.4�՝��WĦD�BzDm���5�֗�.�k�����z�e�� Ɲ튌)(2����5�#=@���S���hZ0C�O2VO#�n���K;�T����\�r�޼��w�rq���Ѭ��e�D[�+�ڶ����qO"M�-<�}���L���]��ҷٗ�SH��^��ČG�2�	�+[��H���7���2��;���S�mn���4�͛�O �a����.<���8�~�g����gB���	�׹�N������oR����,L����O��Z�4{��/�%on���3��E��Yږ������:�z� xݼc�Ti���%���JܰR g̚@"=�o0IB�b6l�켖A� �8�z�#L<ՈY�:ѹc�aa��@\˨�V�{m���n#V��x��>���<K��au�h����d�gu�;u����8߆y^�"��@�`���T�1;wI�/Ok���B�Dܐ�����_F�z�!M.��u��K���r�%��OV�Ն�*���	^��~�sbp��&Ӊ�i�B^Se�}�q ������[���81�ǘ�DM�"�D�w��Sp���G��D��D�����)��4�T�����::2z��� �1/yN��1i���3�1��!�!�?"񗈤��}8o�5����5(1H�(��f�����K�:���r�W%��TWDۋG�(��^g��º95�dro�N�Ж
�
��D����!_语z�X~�F�p"�^�h4;z"�&52I��������F#%[ \��Ng&uY�u	3��UR������j�Cʴ����kJ���5�Zn�W���O��T\w�B~s[��r��h�&l���U0�ъ���������u=����(�W����FVrp���o��M�f�-��{_�:/�K*	��	׺�l��&C灧�������}�����*���j*�uը��ΟF��1�_0li������O��2B���U�e�St|��_�m�+��;/�N���L�X0���U{�ét�V�Kx��,|��/Q���W������NiV���)��;�TV$&X�q_gʗ��Hʝ�~���{68/'�^��������RC~���p�LnE�����bt�%���qF*Ӎ��Z�EK'�7�\<-ֻ@��ef(vu��ZYmyB�'_���Ǵ�3C�n�S�O��J�H�g�B4����,�����n��ު҉���[� �=2�&�mU��}�����_%�)��	��U�;����3�qY��d�OUg*�?:o�\S��w*9�Zx~ �q3������%��r�if�W�x��*o���R��	!���)7�/�R����Z�vJ�az��a��V���H��A�\�~��Y��vإ!<ĳ_wΡN%f�W2�>�2����P8���`��o0�'a��_3f�P�h:W�6�	�(�k�2v@5�?�4��pd�!���X�����VB�̡���&U��Eդ�(2S�?�McPi�U�2����5;|���&�-�P�њ����+�����4E\������//	o�+�Ӕ7-xj ��_B�*��f�/�;�yd"y�S���Ā������1�q�ܚ<<��Z]ɧJNm��ޯG��9�1 �I��i���U����y+���Y�j�;����307MU����#�(юYK�����vO�h�x�S!񥘘��~��WGK����>
��$���m%�JB�҅x9��f�g�%�iz���8��-���b���fi�����u˯'Ȇ�/7=�ߤG��i��؊I���6��ϴ]jiӸ�s�_�ߌ�Q+��<3���8sO��ȧ�ZR�7\���q�c��*q���sZ�����G�_O!����5~�z�Q;)w8y��Hd��O�o� ��9�S��&�v�`^�� ���q���	�#�m淪��[�>�4ɼ�(�$PwA���� &�<H���rƌK���$� ��.zJ�C�G�m�߿/�3S&�o����^Xs�>�t�k#�}V/�\n5����X�蛺4��)���+�:�6���������¢':7����蝈W&������H��ԒK�E��R������ϻ�8��\W_�;Ж?�������;��[�B�ԩ�)�Z���R#_�g(��dgg����S·"�O�i��vE���o�����!1�1 ����k�_#����{)w��-!W^J� \�#��#�EEýK��i�=��/]���xxh������i����[`糼�^�o�0�LMIe��Q���G"��ej�I�:��j�$�]ۓ���QQ9~\�i���8,6q����GDD�p@�Ѯ�Vz���сJ�c't�U�ȫ�Ȋ���ݽ�|�U�ik�x�u��]XEj����&�ʡ!���P5���p��+R���ے��(�e�Z4�@c��.���D~e�q�#պ��N��>!���n-�șH��<:�C�rr��� Ä���_�E��'�L22��<�>>>Z�� �A�a�X~�b�S~J��z�~�E��L��-��&V{�Aȧ&����Ԅ�W�����.���_��4d���zx�ė�i�ɬE$�D�듹yմ��x�z"惤
�4 =dm'Iihjj�^��L"���T���nH���{%a�T`9�O�R��7Z^u=�U�+db��C
����A��6NJ��=����)4,,J;�}�[yn�۾���p��U%^�Hq��CPV������OR$��mR����o��`���JC��-�H�u�B+F��Ç6��ꁷ=x� �,u@�L������ᝃ%�vmc����c���O%8t���������^?�����کS��[>
y�F��25���hW�ҁ�&
�^��lfC@Ǐ���W��;�|H��ڝ1Q|V?ʳ�q����9^899���Q�U��}�����2��3���v�^~(����&���j���v��ỒWJ�l���)�cv��L�>���H(.X}$w8�������`"$�B��#w@(��k>�cZw-��"k�����bm�%h]�E��)����ۿ�ل+�У��ī��-4����5I�Y��tx�+^'ܔԜ�4S%4�5
����l���U-i| �L�����ӻ��[�|0�	���c����\v���ml������3N�_��Tg�H�UY=����4E*��������i{.^FZzom�dHYY켃k�<��v*�~F8m�W�9�4���1��o%9AϿ/��z�Ds8g��,<���z���4�A*�v�!P��}A�!2�Ǥ�`)s>�7�����W/N�ʥ�:��`�5Oԇ��ntGC������^����T�������C�����R/�@�o&��k�B��7
��D�7��[�tᲄ�)䬧�|�����7^5���Q��L�ʕ+�==��TL>0Og��+5�6B����̺���3��.M�ូk��ϯe	?��9O�o�f�7��j�MҎI��sc!��ă�+���/�<9�~�5�+y�ٝO��3�[;ᮊ٘�j6��~�o����W-ws-��E� v?�[e�|���B~:�~8,��*mM2���j��Cg�(\��H?i�C�v\�+
�#���xEnX /@���-����W]Ԧ������ˊg4����?đ]��=�{+7:��z/�Fr��3�>��@m�����ſ��E�eu�9^4��l���V'��s,[i@ἆ��@������"�B��?<||��fR	2��+[���Ow �pRj��w0_�m+�vu�-+�i�2W������ye�z��g��Ď�I��KO~���a��WJ�yp��Ԩo�Y1��`��%2��Ǿߴs�=�>(�"�	���o��ci ށ;!m�.�J��e1�oAߪh��0������a)�.�}���I|`�(X��8��EO���&�0zéVׄs����gϞ�
>Ua>�g���;���VU�����M��BӃ�!D���7wj-�����9�K[Թ;�U^�	+� _�q�X�AX���\Y�mydW���o<ԏ�>�}�z�jk����-�!�6
5$�ғ�T�1�8����"��pE��Ґ�`��eW�W����ŋ]*�5Ր��iqB�T�2��=���f��iiJ���z����&#���/���[��t�8��M��h���#4����Bv1�py�85�����j�Qe�ѹ���t��FE6q��^%S#����56==���S!��M]ş�Պ)ȝ0�k�B�Wͥi��2�u�`J�篢���w�J0S0�Ƙ8]�gnT"a2vy���>�q�{u��f� 0�|Z�ݠ�k���0�R]أå����������N�i�c] �02�	o�./���q�i���ʒa��4悙J
�Sh{�b�l�Tr�5�����dIř�W]�����bk�@i��4_͵��+|�{_�bֿ�ߑ� ��jqj��[Q�K+s��AE�M,�E���Gj#\<����0���dM��ORV�bJndE[U�����<z�h�A�/@&�~B�[Va�X�>�n�mE	�����:w� ����d����:.��C�K�:t���K0�����3k*I������Q$��󱀹<���V���R٥sm_)Xl<���QU��^Ԏ�� R^�,g�[���9���,�J�YU#�b���I�dA�;k؜UDh���F����<3�<��6�;�G���n��$`F11�**��d9�%랼#��X4���f�;��86��4�IE�A�to�����k��"�4�	�E#X&S �T��鈂�j�����j��h���¹6����� ��	�B�.O�-�DpܕY淼�/�����߅�' o���h!�A�|������O����m�h����v���1�l�I�72�m�ւr��� ���A�4q�vg���/e��?@�k,�ȵӻ�����A���3Q�w�Ų��	A����3�{yL�5zE�������rT�����/Y�}>��fZ	����\bW��6ߦ��ʷݎ&˙({Ǒ�H)�>�'@|6����a��E���Ϲ�X|�AW�m`n[���;��Ż̶��|��S�Ar;�Sr�
coǼo����щ��]X����og)ͦ-�8a��O
҈ޫ��g�����|eN�K��%��ǽsg��P3uB�����V'H3uqg��&.� S������P�b��%�M(�P�#R:��m�"��j�I�<WU���d�WWpŃ�-���ϗ��r�\ANU�Gw'M֦����}�c�O w1+A�m{��ܨ�dNz��D��D;j�|�?�����$/:��4�d���������QN�ϴ���Dp�FJL̆mJ��׃~�����5�ة�RN���
����A��j�F���A�e�epϘ5�H{!����]�����"�&z!��#�1�/��ѲL����k}�F����KJ��'�K�c.,�\ ��'X��>@|�Jy-P����q��BG?���(\�j+o)��,�㥩G�LL���qI���1���t�9B�%�Js55c���V�<K�R��H�"o��E��B��zsZG �7r=P��~Y5d�eU�Ĩ���G!�i��P�J9;�7-^.	K�Vݲ���g���[=A+v����|ױ�A�7�o
K<iw����:'''@����4+%����U�h�
�n�T�?O:)��U�-�}XT�Ջ���4i�_�}�k�$M���2J���i~�KX��Ț��$Kޯ�$�H��t��+[�"��O���r�xaԾ�����M� �h�H�'�,KF}�Ň�|��kj��+F�í\oV��+���g��8��(W[9.w�^�5�Dݝ|�ar�y�}M���Fg�E��C��ے�S��.�����ch٬dNNN~@h"{�ы�؃!���e%��_++}��$`���i�J&��t���.�4���_X����vZNR�>y1�iL�!T$^w�'��S���\	u��ŉ�!ϘZtG�4b����Ȉ9�;Ӥ���Ғ�J�w� ed�y���a��9=zd2���ZZ�6KԠ�H�{#�I���T?98.)D�����J�s��sj�����{��.Ȋ�W*�.w,����/���A����B���͜Mjƃx�*M�F�4�.���냺vtl�@�'IY�B��
fw�u�neC�X�:V��wv1���쵻������G9��W=A�M��q��-F�N4��������Y�ң��VSID�)@v��}�+x��F�}��=Jfe�1�.�3��,�^�tu��#��w~R`�W�WAAA����Š�ڬ�� �R�vQ�]	T����6K�Ɉ�-T�$/��<�]�Z�ዬn��IY�?2�����!B��e����<��RDc}��0�)���볁	����>͔H�z����݈׋u������n�(T:q��C4�uh�:�CʩM�u���\��.����g��"��U�!(�����Vۣ��0u�L��Or��Ԡ����~(��E�]��>?�i_��r�k�w_����(F�.6�t����'��(k�X|�o��꣹��A/d1��b��qMh�԰�ǡ�
�\��#N_�?չCR� �E~s�2U��"wl���E�+�_��Nl{�����s(��<:���2W��l����<�rW)�8���D+V��*����Y�� ����v;!1:�0a}�؀�X�|��U{��n��k�j��XYN�p�oO�.��EZ����]�B�ռ���uv��&�3d�5��+�����\��{��*�WEn?V���d��k�8x/U��@r���>Wo��@�ӊ=!"�ǫ���o�"/��(ned���7.766�&5]6�d~X����Y�ߗ/���m���c"9o��d��"�1(�A4�= 2� "E~m����ņ2��AYM�OX!�u����Hƹ��e�Ӈ��V�q��7�1�m��W�hD�+��B�=tas	����Z+��l\D>��-#�=o���*�0jݏ�W���_�]nr#��RQbce�c���Y ���\�:�eu�ۄ���?$ٹ��?��w�Q�0K^�L,&�e���%�n&�7�&����f|X|/��I�����1�sf�x�?�v�Ӈ�m	�e����~���@�/���$���Cm�6�G3��Q5Z�n��� c���������F��V)�Ŏ��Ģ�����9��bE"���k�j&�w��cO�K�1��W�'�N�}HSUw��I��|�%z"ᬱ���_:���u$U�Å;�(V�~�Nh;l�X��Ԑ��P�F�YxΉ���S��.~��*��	Ct�8�2��s�X.j��:�^��2E:aO���R����a�T��Lw'|�"�l�i���gɵ�x��'ѣ�6��FW͜qd�F�i��������x"2�5+Wh�u���Be����I�t����9�VkjMt'��V�`�(�@ݻ��#D�:�C	�4�
�:���=4�N$T�>;�;	O�����)0�>r�����+B�!�ETz�gS5����)/$P	��&��d�;.?�;�B�� �^�_˲anL��)R{�[,�+5��g�..
wSn}w5F����9�:���u�q�%��SV��Yw� �,b1P0���r%7�&�I��5F�uZ\W�����6u���3���4+�76��,�p��O�C�H�x�V��[�>0?sz�Ze8� S�l�jh�v�@"U�Xw�����S�Q����g{a=/�}���É��R���=Δ�/\�g>�`�s����Y �_���.���氂>L�ý�r|~O������d����Uo���]�+E`��E��@oյ��gJ�@��F��g��!�BWz��L��m:�6�~�I���
q�H�.]���y�ń��v���N�����y�� ���/L�0}`� qD%z��,�r|RG�\pĖ7���yN��L��˴J�T�ӝ���)�o^S_F�j6�����$�OƎ�B�~$��E����a2";��T˓�,�-��I�Gx�b���i��1U[�d@~*��Ŷ�wM��gU"�o
����T%�O���F$���	������y����'���e�|
^�߱@������k0/x#<�g�}�O;!����3���e�0r�I-"���/��Ί�3�>M�֌��>��r�,�;E���O�^� J��!�m�mï��Ὧi���䊹���W����RԽ�r���/�%��^�d���v���K4�w�n���Ga�wX��dH,Tt=u��O-_Uץ�����5v�l�.ߐ��X�u#{UF�Y��1t��'럯���:�T��ax6Y����!��Q~�`�	�1�٣>�m�Ŝ���j{;>�
Ψ(�;g�Q���t��D�^"n�2�V�}��1 ��Y��VU��a�yNJ��(ލ7��V���5`o�����_Ƚ��Ӻ Ü�rk�0f���Mp�ծ��U��2 ���jK�+?|HIo�21�G`� �5��}�Ŀ(J~1��I�m����V��j7g��rY�|2�M�s4E/����#�/���8&�4�h�|�xV	;0<�e��4t^H#����Ǥ�)zƫ�ٹ'Rˎ��o��!D�T�����_y��S��&^ܶ#д�%�꛻��7;^�`�V�z0Vy9^�6�uou�rj�]"�(�8�V�V؇�1��������}!�s2l$�,���ů�x���}%q%�zl���*�qg�>vr&�i��[��5���_|ഉ1��U��&��ZϠ��� :2U_?��� -���	N�{���ݯ>��?���'��~Ǫ��'���A����E+S�ޑ��#�+�)0{yJ�n��%z����8�����x@�p+��ƿ˹\����8p쎎6��^4�F'�w�cO9Į^�cr�%J����^�~��vz.{:��f��9�St�J
���#Le�G��H�6z=n1��o�`W��+o�g��"�<���F�[��;:?U�� �˒�|��SRxv�y�Ԭl\R�AJj���nN���(rPG`ަ4��p�ʤ0h0��px�6��§�`r�u�����mv�N=����O~�)r���e,����.a�����O�/���W����m�@��3K�W]-١»�$��ړ��$r�nm��B<��k���'f�إ&���jx`&�_�R	݅ ��٬`�p�C?��=T�=*��$��.Fk�"��#
tJso�?9�j�y~\��YX>mR�i(�ab�A��� �~�����C��9,\�t�)���>+bƺ�F0R��$���+q �����Ҡ�!
��6U��i���vI��Cv,L�RlU�EK���X�e�o_A�~�>6�ŏH �Ib(qTrI�ɶ�FX��IR�\�u�|�x�ͥɁj�1�-�a����h:��������,k��AP!TwUP�"]QP@Z��J��KG�zD� A:�C�	=@(�|��Ͻ�����������9s�甙9S҄�{�|e�A %v��=3'<�9U�ԒN|ќ�nM��XbہK�ڃ��,�ӑ
�w<7�6�׮�K�~��-��g�v�Ս]0fgVQ.��{U��yt.� � �w�v�h7u��R�9�?!�:M�=Q]k���ء��;��� �(�� LYP%k�|g=>J�ܳ�S�0�a��8>���p.��=�õ�#ůY����Z%6�F�Y#΂�Ne����<����u��S��L�nt����5�D}݂Șm��Ր��x�{a�r�ܿ�V�x�ᖅ/�v�J�]����h���bz{�Ҿ��E����
o/i��������H���k�;�}Иn�Z�oN�����8Y6��9u��=�W��c�ly�ӎ<ǀr���3~0:^{��Pm���g��=����Q^XF�.W�����~��ǈk�+�aG�8֒}hkMT��s�w_�MI��m�VaQ)z+x7�Oo��Pl��q�O��W��6�ї�)|V����a=�l�Pva
��L�-q�#��)�{R0\�@y�Yb�0x�u�E�/�i�#i�|�k�b��tJI%�RC�?w�^Xn8��|*������'�-�?�e�9<�fR$4�V����<������y �Q�%@�q�Y�'�k�d�W64[<����ɡM�eȺ|�r�E��V��W>%e���y�:yczcF4�����.j}������n�31}5�,�X�d#���
�!P���+o����ہt_:音=�]68E��ˌ()�������<Fw�^�8.o�5��:7ݙ������K���LuV�_@x�����{��M��aj��⮶��m�2_lG]�)
�(��	�ˆ�alR��#r8�:S��%)?:s Ko|�60�m�۟-��w$��b�#:K�M�MIzs���BӡBߵ���=p?�N��`����� ���8H��j������~$IX�n�\<[���}U)CX�'��e}4T�Ua$��@��I��mo�M?�W�Ś����Wjn6'������IԄ��FX���f2�vY��>z=-C�ֿ�hH�I���;���P�:� ���n��Y���ys���7cx���t�E?/H<	�P=_M$)bR�����HC_J#wZX���SPJ㨚�a�v�!\t�"C�ѩ`�t���3.S��+��!�}1ݻ�m������lA�g����O��*Y��Vj.��M�I���P��R�;�hv��a�f���qC@9[�3����?_�����)�O�B���2�-�b{��V:��P�g��a������� 	��"��7�F�ﵣ%���_��%-�</�s��X�әU����K �����8���A�J�Ջ%6j��T�R;�]���}�겂�<*��[��I��sk�U 2z��v�7G�q%H;��(	V��K:}zEtRoo��8y�;�Bi*�(I��g���w��/�]��~Bۖ�f�ҞD���G0=�&�[�.)u�"�.c� ^�����$�i��@j�M���)_KP0�gl\g���iEԶ���<��9q�w�R����'߶;��k�bt>T�y�|"Q��8�B��E]���9f�ze���4��V�)�#V�Ћa}b����(��.?|b����A�ɬ��ԑ�%r�
�(�lUGR/�E9��.ٚ��y��`LdfNE�`��>��RV�>�U�M�p��M�X<�j �Y�)���6���o�&�0#J��F�MS�eE��K����4.�g|"099y���%[I�RY1";u�'�}ݬOW��nʤ#��})6���,��V���>S�K.�k��Зn��􆧚q^��.sX�qFb��p��~L9R��3H����k|�m�<�N҇j�jSw�l��Y�:��-!�gn�����m��E��_hL�Q?Nv,�k�M�!���]��=JT�w�?~����~�Ѝ�dy��*_�����2��v��-t���Cw���V>��R�^�a(VD�4�Z��]H`@23�p=�v\I��
�._��JܸW���γ)�����i���b\cLL�P�m�����=9��X�
��E6v[me<)M@J�^��Q\�ѣ� ��~~���ZL��5�؂N�ϘN����-+<�b����l̢B�{�K�;)ʊ����|�ϗ�{{{ێr�!�h�u~t��1�.�9̖p�y�ISt�)y�Ҥ�ECc#2&��C�10��{�j�ڠ��_AW���rx�0~-PIF�L-ʊ���~ඨizL�J��O��߄y�e�~�|�ZDv��*�%�:n�Z=v�.�-Mb��!6=�ĥ��g�2��vٕ��v�����Z�U��T�E��^��gWl�{�J-�s�����"�Ss�,����ﰌ��mD��aiR{�����N�T���-$xת K��z�R�Я�_O�×	����XI��HF�y�=)Ob�
Q��UJy��<�*���G�N�K����Y����j7!�R����V��0�;v�x�R���T [�`���d.	���P�fj��]�c߭��?��,V���������,g�lҚ�(���˲
1�mé@)�'�:/tf��z��ݼ�������̃�qq+Þ���������(���j����{
R1s|m+��a� :�<f�Nuܮ����!�Df�"8���W���~'��a� 6�ˇ����~�+��B5�Y�u�nP��ľ���N���(����OjM�I�9G�@ny���&�`
)�j6N� bj���t�]|u�E�L~+M?�l�%'w�b�'@SRT̗� (�h����*���������;2 `����zj� * d�v�i11��:�u������'��6%%'�*�d��\X�Y)�S��V���~�\3���"���@0� ��mT�d)����;G��TTT�f{r�w(�>�<6���c�$�e-4�!��e�j�u����u�]�����Ri�-�����1---�E˿1��z!4�mj�>'��6� w�yH:|] B ��(����4��~'��;� %�u�
�	;�"�1򷳧�[�s
��iy{���B�ҕo�k-PY!O#��l �-H�2�ӵS�S@4q��an�KP%����2N� �̚��Ó!��7��Eށg]��3՜�Iq~υ�~ ��	X,�y�Ɨ���@����]v#�������_��� �}��J�j+z�}ez�ʂN�a/�$$�iX}�O�w����d�Ӣ�dM����r �Gc8��ٯ!��.�����_��	�Ċk<�Hŀ�7���5�%P��,�ɒ�~��nw�y,GQ�^f����ߎw1-mhԎ]�z��`@R*�Ĳ]�E�	8z�x�I�w��X�S���o�j�:�gg�n��o���
�6,�ˉ#�ހNr�~�E ����t�t�����U������\��"xSy���� ��q8������v7�����I�A
P�/��-���N�ϱƗ�rp�q ���#K� U�������m��{<d�o�h� ݪܴ�yW��~a�:d}> ��v��@p�5yZwY]��1�m44{�l��a���i�D
��ޞ����iu�҂���֌1�;��-d�
f��t��n�o�W��ٞ���)�)j��$��{ZZV����Q����Q�ee��s�v����ͽMH���אZ)0��s;�L�4��&�ᄄ7D��9�IK�����(Ah�7��HڏݎE8����}�^33775������	��V�����t�?���n��.J��`�1����� ��m(�ܞ������FUM(�{�!�x'KP�����k�#��~�T<��Ú6��F�d���~��	ĊW1*���Ħ���X(�.�HC)�E��c����\��8M��A5�w��FgO=��dTP��6m�2���/(n4]�����LI鴨	�U��&�]BA9��ʏ:^�A�O������/�Q�8b+�vnJ��K�2���������2�Sɡ��8�BP ��2�#0� /��h��j��>���SIzJe��՘fh����/���اW��z�"���N�+��?C�+�m��b�9 ED7�G�H\��(�6F��7�ܦ�����v�C�Pi��|�d s-��a�r�E�C�\��ֻO]�����/d���n<謥���*����K�$e����Z��%\���6AqǾq�G!t�!��yw�	�|�Wfd�S�<��9q+4�N���f�MFW�G�:�?�T�}k��u{�4�8'��� ����J�&
&�=ؕ`��9yy���S�n@A����G�Sz���8G�Yo�ԫf�h��@��h�kV=��_��UH�'��r�H��I�s<k�lKb�:��	��(V��CG��b� ������k5X��J9�?����JA� �*~@U��0.{�0{4�}�h2)Z+��t�ڻ�C��淎�yQ�2���p5p#��h�����ڞ�.�Az��
�#$��j�`ٮ�DC�+�޲�v9%�<�H��S���Cϡ��8-��Ժ�U2�nh���e��
+�P�9 �@�߃Hw ��{�@�����d�׾s gM��R @&� �A�nfvncc���!�)�]�����B����xf�Ũ)T#nGq��)�:zX�[Q��η��s���x^FFF� <�B�y�j�uc��^�����`�ߏ��u�W�X�S#E}��4G�>4feʧ]'=�����fv��q���2 �����r:�
�������@��2#�p9�W��C��@�wx�⏸ot�B9�ͣ��}�[�P����d�V?($1�Z��ʖR����p�ii��ܦ�2�g:��`�F,�ɪr�O�Rq��7�Z����9;(*� �5�-]ޑP��Pf��>"Pu�-4""BY [������8�TB���Y4��|h�֮���ܮ	��Šѭ�:z�ijiힽ���bfީ�mM���+�r��kK��T��A�y����J��zKo�R}�^^.��]�NS���O������F��*���f(�� ,��9f׿%<� �VXq��2.�M��^%F�-F�k��q� ܍K�t|���S���q=#ʉ5e����h�*����p�w�d[�-B�$	<���w�j��:�m_]cȟ�4uɱM1vhҘ:Ek������L5N��8�CqL뾄�ⓢ--�X%�`׻/ْ.���,�����S���`�ssj5���T3h����@_d��r1��'���/Z���Ũ�S��ܵ>��r������D3��]ŭd�����rp�n�S����"bg�h�U8ݮ�͒` �*/kl7 �_���7ٿ8N�����H|��:��Y��<p�E�h��Q�}���<�)O)����f���/��W�rpqz��芦|�f ��M�_�e#�s���0=p9�ec�4�<��H��}	C��nv�ck�@��;��8��- ����Ui: 3�|�hi5cLķuw�̓G�@xe��9 N3�H�.]���/���Y�?�H� ��p��Z�IEx�Z�0-?~��������a���i��1�?�D��WK�b�+7
[]{�f`N�����r2e��!�/��P�w�Ö'v8�5}[>tmt�V�i�ss(�x�N�|u���/�"5����#�u�N%��;���Ϝ����`iD;?�t�d������Rk{&U"����{���TP�k��[<����^������D����lJ����'Ų�Ϋ$�y
�U|�H�M���.V_�,B��.[H�s��X�l����g�6�����q�'��`aM���?U��ۊk߮<U7^ih�'�Ғ�0�p��_=R�kz���x�"��Qtn���ץ� r!̟M�[ګ�2�Cc����"z��������W�/ˌ"4o�ꗾ��]��&���k6겭�}�@��,�@��Sd�4��8�����m��zM�Ym2u����9����>��������Wer�Z�I�T��/�V�f��7i�C�-qdKf(m�j��0wf>���-�sಜQ)]w�.�Ħ����t{5�k_����Z��R��;�8�j{{Q�W}���a���ո����&{ٛ�`u>j��R��$����FX�����B�\9!O�?GW�V�g$�Ό%�oW�7�M����V&�_���P��A�窹�KWsf���K֤�p{�-�$
I��7����Pd��_�g^�J�\c���|ܒ��#�	'���+�B�0�}z\�*(D�m���nSg*�KǿMn�h��4t�����Z��yL>U����+�1�zx��uS�ZQ�!���Bq25�@!��v�>Fjj�� �5|L��mT���J�[O�' diҤxQN��\<�̙��E�G��q��������V�Ul���/y-�3���(Mk�Lq�M�G��yjx�s4�D�J���P^���@&�ңfF�މ~�s�����sJ�ǂ�mmtL��#�褠K�H���W�=����e�]�&$W_�����R&�ۑ���%�q�N(@z;&�`�3�[��n�3>��I���An�����VBԭ���S�#���j���}y�2���Ѭ}R�@;-_L��/���K�סg���{R&�?����DFW�p�����-r�E�5N7��'����\F�	���~cܒ妮�H:��k��s?�}�+1�<Y`��*�[��^�?0�X~i۲���)��>�]��������7�%h��r@��d����jbέΥ+G��[�o�_ q]���Cȁ�������!�QZ�pi�������Դe�Կ;u�+3�Wዑ}��ܥ�B�p����fmog��d��|���v���c!W�
��[��ǣ�"�Cy��ff�)������h����J�ϥ�#�[R)1)lpq8Gu)s-9v4 Y_��l�xj>p�Le�1���Ӽ(���EֆS�&��Xڵ�B(��kے<�e�cM�cw�X=<�5�S첤��Ի�bn�����O���l�)\���0ԨR�LگC���"�/) O�p_-���|�.aHnً]4�a�{�7x�D	�xb�܌���� �)��R��d�I궃R�B	��>PF��Z_^|3���������'*W�8e�h2�@����F�����te��/�{�}Ie�4eU�v��mll,3.��]fI֔�R�b\>ݭ��$x%ELJ��[-læ��+�HI�-���34�f����=S��Q5�QS��twN�sc���~tl�������7�N��4����N�u4���z������T�����^����;ȁM�`wc�k�m-�mx�&1�����Q����35����2���b���JA�� Cp[[*�T;|��4py;j_l�o}��b��B���e'�������)ug(y�l|o�[uOᩀ�[c,�rB�kn�/�O��i����%�G%j1�}������������L�%]�!9WB����5?_W͛���}ɺ���R2�;7����P�©�h��R��9�b����^ܤS��@�A��8�fi<,]����XNv�Y𝿐O)������P�	nA��LW��[�uF��ud��W����\p�"��� �G.'\�,&)3�ť�U��	O�隭�W3W|��!��q'�SiZj�0�d.��(Q@�J=X�+��lP���5�
\�u�#��ta�Tfwi(/��R����v�K8�b`�9�@�_��Y��z����E��������7�ٝ9Z=�m�bśT��#k�7��3V��XY}Y*�j,e�Rڏ�plC�����]����>���z���Pk�x��t::��b�ht�\_Q]	!���d��{Q^�����[O|^D��`����ތ��\<L�/��c�L�Zx���T5K��+#����Yg5�ð�F�&��=��.��%����וڛDb��]���9��6A!k[�KF�������aכc��[�q}��	=j��E"��aN˼+����y�D^��+J:��D"
��F6f�A�1�2��E�Ǻ%0`���FT�/��P&�]g�F-F
���fL+����}�����J���)��6B��ySݞ��,���*�0D�E�uԈ�r293���m)R���̠�3���>E}�H�N4ǘZY	w�����30C?����%�b��������i`���	;M~s�ŭ�g�Z�ϟ��4��Ͻ�_tp.ɿ���'���6vI�n��<�+��v�ߝ`��;�+�A�l�纇?�f�N	�K1+���;���q�^cZB�= ��k��Qʂ5*F�!km6>�t�\�Zy�6	���`��۾�����繐R��W&A��VT��2��w��c��b�2�m����ks#��wV��x�M��`�'Rja8e�@�W�����Ny�-xY����y8�,!�L��uj�8,'��uL��B>�^�Ⱥ�!�/�d��?����Ny�0,�5P���@��`P�������> }�=iǌ�uIS$RP�~Q�n�G��s$'�n<pxOE��R�$7�h�8��4Z5CV�Sjҍ����.���i��^�3�~�k�6k����Kͷ�y޸��@2WV�|��9�g���$
�s+��_%e��o͚�Te�
_����
�j_�Mzgm�>#"PwCn�=�|r���d���x�8�䳸K�A�=�oXVȊTn.R�(��~�lՙUd�/-��mYl:&Rlҙ�(=�*4H�#Q<�w��J�փVj�7�EQz��%$u=���]���Tn�U��Ў��������Z0���b��[[qLW��b���vB�<0�^��tUx��GX��������4T�@fm�%�)����ׯ7�z]����^}4Z`7�D�q"ı�;���@�q�E�2�p~\?cz3Y���w &��0vJ����EZ�Jy2?����6�}��K�F����Z]K����ʛ��638#�l��/ij7�c�כ�(��
'��V��q��G��t�m�̨���?����b��$Y��9>(�,k�����}>J�e01�/��w�V��3�֧Wߧ���-��;uɖd(�2�I!�N
{;Vq��%i::_#�⸲x�{���~�z]@
^�B��l���� VOB�nm�����l�ş�)�u�W>KG�
��)䭪����n-⤭>���
�B�~�
��#�B��E��A�������cXK����S��Myt�:I���*��|;�Ⱦ�~�P��5o�=3�_�<14���X�j�N�n�fӐ�8[ t�L���_r�3��b\
c�Vb-Z	�1'Q��J�x�d닕�־ZR)��C�u:H��/8 ��2x�Q�5w[�t3O;j���Lc۪�C�3�k��VW�+��C��X���ӂ�����G��F�͊n�O �[�q5��w㽉�%,D�س;�0�"D���S���ovt?�3��şj�e\��_�D�i�Z�#��e�����~��bR�k);�������{ G�!"ͥ��ovQ
h������Y6�	I�{�T��w"(�}ޑ�
I�b��a�[[`��@�����8�|�z�l���>A��XoԌd6'$��R��gx�bNp���[�q�Nh��<��A#��3�,��=��u�^t�yFY��40�S��Sq�렌��E&>�Ĥoԍjiűa"��'���Y�#�^^���uY����0������6�l�%or���y<�!�ln�n�,�gW+�m�n&Y~N�R�b*ێ��|�ہ+�<U��N;��)X!i!���_��Y� �$��&���.J~��n�+���]�ܿ1�cNx9+�D	܉�T���O�8������_��c��b�=����s�9��G1�����֣��JO�����3Z�P}'��Z�S}��cr��䁉�/l�o����t����Α+�mY�R����٧�����,��[�SG��+�R��[y�� l^��.uvypm]�x�A����{�?:���l"@~gI~ga����n�o�p=���*m˸��L*�������B�Y	\A<����8��"��^���\�0�_�8������I<�n��|'�I~k�L?�VQtron�1bK?GzX+��r��ÇP���^�!�ԝg��[��7���C��Ҷh%�ytE��te��qU��v]bRX�d��kv.���y�ܲ�s��cW�E?�</��!����ӊ�;�4G����u��nѼ��͆2��E�5y�N��ݪ��T��]���U5�����<9�CO��I�SYd8��^1��G;b<��zfk�fk��7���fY����F��g��r�zK��愓���+��'�.��,���,����Id����uu������D�(�B*���~FcF5[�h�-aΦHіԔx)���(NS��;�q�D �CS�aY�����;�esVO��L�`a��,�-ϝ;��2�a���a��i�ˆ�Mdӎ1���T��TL�O������9�9<��S�ɒ�降��q(��7������VZ�b��.�����y�= ��-�����bG��Q�6J��F�����L�=���R������X]���#1
5�z36܍���U�ny0�,��Ef� �����P8e6����,z���!A�+j�o>�e��C����B�̚�g��|�@m���^��������xL5ή��A2KN%�G�����d��EE����`�6�Ʈ��ў����z���E��%"�����:	̿�aeBE���E��X��S�b��:����EǱx?z9��P�O�E>�ϩBNƺy(mKN�l�#у����><�w
P�fU����,��[��77��ѯ�${u��)zM�F���Λ�e����U��G֞��=y��'qm�G��j�1|��ݠJ)ʃw��=�[AW���A��TU夂���[�.�eơ�}�zJ9�+mQN�Y�U�ם.e��O&G��ŭ�Q�4Yxܩ���L�V�K1)������I�����,��'8VF/2�!I�z�Y�����;L��`�L)b�D�w!�pH!'?u��'w�ɕ��-ɯ�yI���q�b����W�C�~��6�I���e5��z1��֕gq>���Ք�:�d$�7S��}s��2b��u�F�p=J���md{�LA �`7ZI�<(��� �H(z�E��j�����[dWQ�ѣ��$`�0NS)@��Z��`�ԕ�u{�6|.�ol�LI��JM"��-]�_�m�'����	���n[d `@8-�*����-���`ƶ6�pf��"`0�������?�7��є�sQ!y�+��KeOi�lr4��cX�3#���Kfs�j�tė��ڃ���z���&pO�r%�}�.���󐎽o"��<<P!qJx���[z�RS�^�U.f�'</f�oq�56Gu���\�R�nvN���_�7��a�q�������\��b�ݳ��L^9���ᩇ��~x���!�W�ttI\��?�z��6��/tO��TM�;���G�6�Y�ҳ�9
��D��O�����@��_	39�����%���%��7	V�?�_ �?��$����T�'�bމ@���%��7V��̂��(��������@��������+t}�IHHD��:�}�������:��0���:dc� ^����A[�g{C�+�n�T�����5�L8��r^m��*��.�DcV�OL/�K?'�z�l�?�3�yl�������5�����ݠ}����t����x��H�[+�*B�bT��ߑ�_t��N
	B\Sh��g)"�)����Z>Wd�4f���>�m�j����318zd'B�%��ܞ���W��-�vE�^�m����)���ĵ�L,�Z�30�W���U����[7����������P����е?E�Q�\q�_�ɑ#�j4�W 3��@����ϴ����9�Uֆc9e� ��;ۄO��c��v}�����Q���o���,kY�M>	?��`%;��y
P?��gg��x���(���7gnK7�t!�� l��J�=˔�VM׉�6�^�M�ߤcd�7���=�7����|GHdJf�p4)p���]�* �y'�V�'i������URQǎ+�U(�Wg���A[������9�}��y�v�c��g/��!����o>�m��㧍�$�k�kM�'n�m+l`&�E�=�e���o�1a�hi�
;��,��K�m�߷��+�ݤ-�P�_Q�\���W�AX�.������H46�x �{G�6�#����l��\��kS�~�[�� �m�q4�%��+��$����,ƙ�[�+�WW�=���g�-�r��A{�W�W��_ �24��ĹW:�����}�&赯�݊o�f��u�{����0��j�l���c�V�m�v�����ـ�7�e��B{{{�~����#(�l�o9x����ݰ����{FK����j_�҉�f�s���j�V!�J�wre��reӗt��f��3t���D|L���4����/�
��V���mJp GPh�� �y�����b���G�����cM�i�=� ,�`υ�F�hj"�B��?�V�ޮ�H��Č����Ə�)q�.��p�.�S?a~m_�S��\2���lZ".�/��=~�͗����9!�n��8œ��u��1ѯ��M,.�G���l�Udm�?��{�����oj���Ɔ�0aV��]aV�V��g�)�s#/1t��DG�yQ���`���F���Ƃ�y�� �֯�+�W�j��r>���@D�R�2���c�j�{�x��V��/�4T�bu��6l�JT�8��Bx�D<�F����1237?�^	���;�>��z`>�j�	�δY�4����5�m!Ci1��F�yЇ��V{�����6����p"�c/e}I����n�G��bݏ�V���z[ܯ�'�9l��7G��:r@�6�|���̇���\�&.�k�Q!_���rsm���؞VFdwyQ�lA'�qK��*�cam4�p2a����G��6���'M�ϙ���?:D�*n��g���ŗ��Ro��X_^
����xnO��Z�-"S��#��׬�r�zT���X�d�$�x�}�����KoS�,dm�����D�x��t�┬����D���1�7YK��GP�V ;�����vu�8v���$W�4b�� ���D�|�ul ��JN��4�͝�%��Vs��p�n���mZ��7I��ˀ��.�&̺��W���m��H�X���J\c9�0vH�MM���r����\���1ă��&�ܢ���ty,T}����ܥy�CWt�M�l{{�z0�zp¤!��u��CĤ�X>��b�`n<=�AB�ki�5}6�=u~�V�7�"�t�m�p����[���=e����&og�V��/�p�ז�3b��(��X�E�e�6�Jǔh��m|.hXr:U�HPml^�"n�B��I����X�`��N&6���,��_�޴�A����a�4r�.4�/���>��%�����L�|��5#ٺԶ��oG�d�EM��U{��������=&�?�y����/C1�ĿԶl�X��FY-�?��ŞjD���J.�=��g!��i4p�q�%堪�\�k�]b�#C�_��t鷓�>���*q'{����%#��^�j�p�ޞH	<z�/�8.����l9�'_�Q5��Q2l~ظ�ͰMS�Q����u�������F��C�6�������܇U� a=��O��͖Pf=fդY�>}?+C|�p��X��Y|�x����7bw�ׯw��K�.1���'�vUt�I��bTcUA���(�Bv�,��3Y]b���>Ԍ�x��Q���v]�a_}�q�p����U{��q|�ك��ǸMu.we�/�浜72̵��2k�'�&,y���v4��Z7De*�����b㔸�Ƹ%;lBq�P��ٵ�N#�O1K]/��vA<�)`<���G�L�8g
`oQ�:�?�p~�Qcx������Rx��M�cڪ��~��u2�y�O�|؝;� ���wF�u��<]�������s�7V2���a`e��U LL,6۸#��S�SSSV}��+�Y@���{p����ߛ
"u
��R����_��qȼ�^y3Qh��
�HNE'�w�þa��x7�R�B+%�bu1)��O8������b6��۞[�0��z)u�bOO����gb��HM�o�;����U4^%���8l0ף�g?��x�:��1K-�|{r�e)	�+op=n,	�yV�(�*�֍��Y�r���sz��7��Y��A�57����>�o�D�aм������֙Z^�%l�Ͻ!����t@J/�5s�R��݉]Qy�f!�j��)����G��楀�P�v��AT�c����]F�����*K�V[ .*�դ���'�k��b�~Rғ�Vpb�ˇ��kMV��4���ҿ`��WM��W���Ɵg�k*�]�=��43S�t��!�<f"�K�ؿB�V�7�X����o��6��Z������=D|�:d�%�_ߥ�Bm<c_p����ۚw܁@��3�@��~�ǟ�5��.I���$ޤ�D��R{����r	zx��J�z~���y�nLtKWjZ�Iu�2�G엣��,�E�1@:W�2�e�B�� �TZ���p}�t���I��;gk.��Z'�w��\tqG6�n>4������Y قș������#�1�~|:O�i: �U�c�A�!\���M���.sO��f�}q�&*v�� ���/�5Im��Ffl}�ٚ�_To��ӼR���'������\J�Y76��~�<��m}XʥC{5  ����mԤ�+����]�]�Ƶh�H2W���Pf&�I�g'a���"������-n���M�R��`� {����8�����Y@�Q�O�w.��x�$����7��ЉcK�S���	"�n�_g9C�F,���Aπ��G���0�'K�V���sA]���Pg!���4NG�>5q�L]��H��}�w+��>.Ԭ����xB���^�BW�U� J�U���h �ۆ~GI���8Z��P8�m�ץ�)E��G�ڞ5M�א���ęC�K/t_����Ԡ[��Nj�*�w[�aI^~�@��e�h�=�NMݲ�=�b�JϽ L�Q�3]�$d ����E�v���"��#���R׫�7�Dj� E"�������u)��Bw���Љ9ð1!�;�?��4to�a�����X��	H��]�փ>�µ�50�"�}��E.]9D�&��1Us��n�jІ�D�Xm��7��بǷ��[��7)M���D�Yl�.J?�a�q�ٯ�]H�����J�SV|������	sUe�(w�&N�^��j��1�g����ɪ|�wƛW�7g���i��1>�]��C���O:ޣ�R��*��P;�=&m�rn���0���w�p��#Zi`��.�ׂ�W��S�*�6���u��y2����ET����Ε�5DU�k�.�>��NdAI���wΉ���Q|�`�z������V>��1������M�Xlg�.��F���5#�X�N�H���ȓ��3�d�#�4�16�t�����n��U�����!��S˯Z��P���n
��(�+�߉��f�:�f5�\I���>d�*�Ib���Nׄ�����SY�TA~����0����̢f�l��NH�ӧ���v��H�q���TZ�w(�?�E�o�O,��tXo�ay"��aL"�?���9���!LO.Ht��Y&�|����M}W��p��T>�m{-e��ǥW�Dͯ����:镅C�����x0?���jML&J.7���cU����%���3�i���$_{�M3�M.���ۋ�|q��� MQS���M��x�k1������"ቡ�5~�G@���?8�JCB���6����%�.��A<��$Kh�^���y�ܼ�/��{���~���Cr6���v�w#�q����^瓜:K���]Ľ��	�����qM�sE<�u�?�j�Y�h��E�̷�n��%5�p�YnE^[n��3�����ƺC���O�!��-N������譡��a�f�"w��L�ݥ��,f���a�.����i"�-����l�������EK�ʃH��;u����N>}�F�B� ���jHX~���=y>�n>V���{ay���l,bMϢ�_���7dt��x��26ͧ^0pS 6��5�w:�g�c�(��kn��6)�x���3FFN�F濧����~�����"+�� ��]������e$�k���?��&�1����5Ɵ�:�7�*2����p_��QS���/h����Q��>U�b)�6ݶi�:�4��h��S�Rҕ`����бe���R�	�c6ӏ�z�o��gy���%��R^�+�А���♅�]��Į�.:3*l�H�ם���4��·�|>T���T�+QL]F���q<_}8EV;�]�b+0>ouqq/d+$6~�, �)�`I�@^��޳|�*l��v��d�`_��@\�sl�����WjeR�.���{I�(�%��V��N�BvB�̜c���C�v6���W�y8�C�?���#4����QO���2s)����k>c��Nԣ�%R��;���s���|o�֣��Ӆ�|5���gG!�������^%��*l�S^dɟIg�u���O�G՛#tN�.z��M��8���5��i����ό���y�ȥ�U��,>̀P�7�Ɵ$�[��n�
�0�*OM�5��r��ta���7�rZ��@W� ��Kw�z�DU�g�&�'���v5�Kd�E&= �! �dk��+]a��⏲�W�녇�t4�~���+�3��j�Vr��9�LC���Q�	)t��L����(K��T�w��/�Ԇl:͍sfҹe��E�WK{�BB7����*-���e&��'MԱO�ؚ��x�B��鉲��"�K�k������MK.=��p1���y�=����PH|hr�b,^��Ϲ�w��l�b�f6�<z�Oʽ��қB��$�Df�7�p/�|��s�;U�1���7h^��V4��?K㈿�������N�D�{��)�����_�5���o-_#O��SÕD�c�~hg�䢸�O���J��>��`���|z�� ,G6�iɵ����pa!,���P�LOJU6�������j��!�����&�,Dw�`�N�YE��W���w	�d���'j7oa���0A.�coKl�����b��[^qtc�k�@��LM��'�o���P��	�;���Gl:`����(I�e@)(O�]iB �q�W�>���K%�*�6t�~]��k�ub� ��;�����N|:�침��{�oU����'<q�$�T>�����ys��N�R
!}4��-t���Ѵ�
h�?�e6g��Z���ӫ�g1[���.B�B1��3|UFf#Dڋ�by<�K��B�?�W���3����d�M�����3a�	~�o�!w xh;�na��Ĵ��A�Q���)%�#W�`&Uǿn&�D��������MvN�R�U���G���Ն{��9!!K3�Wϟ��8�~̲{B^`}���j�k�d��>��R��?���y��Y%>Xq���pGy�j��I'S��Cg�*��D�k��=ZP7���L��\�^m��p��UH�%>D����$�������<~���#t,��U������M�	�$�B%�7L�p�5�����J_=pz�� 0����/��iĊ�W�v^R���,�nt+�A�Y����-�%��g���-�x��vt4z����[�~�����Z٘���2 E�*ݴ���o����L3�M�*J�և�ɠ��R�8�9Z���� ����Ak�����P_{Io�^	>�v�p'X�����������]n���m�L]�̤Ȭ�!�(SfJ����1��2���)���2Oq8���1��]�v?���=���Z��z=_�����k�j:\Tأ^/v����uE����R� }G^+il��>ɀ-,��su�nl���R�ŏO;+�[��[ ��D4�������s�8z{-8賡a�/�>���~
x��$?�7
NF�rg�m�B6�=�iz���Ʃ�����眵�KtZ
���:E����O5=�dm'(p]*�H���B����ss�V��E�9��>H�A�H_x���I�s�}�m�Sfqc6��/o����C�p���J�u�����=���/8[�_��-���P`>�iKp���ε"�y���`6!���e|J{z�ʂ��p�ιy~a /!]���7�[�c"e�/6���(���?����Ǩļ$��-��+2DL�u3P�
ޡ�/Q���z@Cu�V�iH��8�P�{X$Tۮ��?uj��^ps��[WDO^*��nN����%��C�gdt�g"��/��xC��E��%��B��S����ŵ�z$C�b����0eu�9��\t<����5�=g2���+�5�/��3��e�9['a5�G9���7�뀩��.ǧ �O��]2�هac���8h<��8��腂-{���.�=6%r�oo*��"�2;�C���E�J���Yl��6
K&�;`�=���f�4�9kE�=��}��>�rO���}�<���	�R�{AD��e%�H\fy"��ۄw�f�i
�E�梔�tv=���~����}�zd�^�i��}<d�5��kg��Q��j�=�{�P���0�6�1��lW� ����BH�3�����f�Z�>���s�%��\	�Ǖ�LOd��ٞ���p�{J|ieI���5p��Ԋג�UU"�:F#�n��쑛��[?��'� X�**�p�O잷m�z�lA�k5�D/
T�/J$�+(�P�J��Zy��'_v�fХg
�cQp�^챙"�^{]��4Z{IDi�t�{�^����uD�v;����K he��B��k�(3��O���}�Xk�[�wZ0�(���[N���t��9����4?WT�x�7��E3��)�tW�_^�$-~/�����U@;B8�����ʵيhx܊����,�kU�������mω��, g~��lf��"Ҹw ���,l�QT
�$z�~��r�.$P^ ����߼��U�C��\��ֿe�0ف��?��d:���&�m�`2hǯ`*�⬿oL�!ꣲ�u����R�ZC�ݲU�v��Ր���@�\b8c�
��F�}�� �2�q"� `gO���$�y�#��y�=����q����:�8g�`�t�.t��B
Ȋ��S��4}�F1���6����HK�ٽ(W��W��c�)����n\�iȗq۬��ת���.�x��g(7���?./=o���b��)�y���R�bL�	�ѡn�۟���kfC�~�'��S#��p+Ng��Õ}���z�I9��?��^��U�2�m���1P���=Z�a�l�	�:��>�Qt_�G����P_��[�Z:��ON���qe��G�p�^ n���\�9R�]Gmi�V�ȯ.+�ߡ�������V��
@ș�w~񫋂�5�����{�G3���c���{���V��/WdB���wVQ����"�h ǭ[Ğ�zY���(�u8S">E(n[fɷ���Gr���B���aZ)H�N+6r�R:"�e�F� �W	u�Q����S�6�V_H�?j�|��{V-(N����(��:�|�\w0��Z}]ۺ�{����#�a��ur���z�	��W��4�7�)�4��B� \j�Wj��7^������J�θ�<�7���x���p���V�>���.?��u�
G�2놧��!��;��C���+�ƕt�3ٝ]���
ؒMk�3�_�M����)pq���Z��E�U�{	ɑ����Ķ)����dm5��h�-Lz_L��b�(���/N+��+f؂V<J����t��u��@/9j�DWg�����%&��D4�w���V����t�1�l����A�ج]���S� C��)���(�bUT0:�?�
@[��+�8���e��3uG��u�6t=�_���N@��^?V2�PI/!�v��0hX���솘��<��>gJ$��h�����eFھ�%!�G�&��R��/嬝�C��O��4/|G#m����i�&�f�D��^o�=�A��ske�c9�Iolǣx���{jq�=���9o��\�����'�,l|%��� �[�@��$y�������L��E[c�L	�;W{Z1䱃H���3DM��i4��1(�G�bhf��
��x��x�� \'s� ���G��Y�D�H5����G���Wq��#���"�#їP_�d����7� �d��X��:�~t���p���E\�ФsxFF}th�$8���7��7�e��:�Yw�� ������f`�&	�˷;`o2OF��X��� -��8�}�$)���O*�H@��HM�Ϙ�J��Ģ�w ��:[f��E�����^�HU�z��0����9B1�S�T�#LLv�{�U�lRT�#$�(7}�u+���C��N�Խ��B�b0]��JC~�M�C޺��t���Ǫ�[�#㵊��ď�3�(����S�ſ��eS`F�hҹ"����e�Ѽp������(
���	W�*1��v�`�gR�X�������?��� z���gT���L?֘��T��m��B۞��v���9G��]읠�5dzFd���`�������͚@[QB�g������A���M�a�#��"!�P@���ܜI��dQ\x�F��.�f�dC�J��P����]��
�m�����������;�.���iq�yQf���15@5[c�rqT�hх˙��J��c���t]����M��w��>���\�-� ����~��n���`���E\�*S *^�6��-���:u�L'X$)�ג����}�K�q�;/���/�
��"<�yzgBbz{�=S�E��itz�[���V1�r�U�2�7�1��:�΋`�P��b9;��[��Q�<�Z^��9M�vu\]�:���W2�]5U�i����t�������	�؃P���)<��`ke�m yF�K�s �_�멿�\�c�t�n����)��vE��??��`�ǵ���ygi<^M����;�~7��)�%���9&��MpI��,ՃH0���gw�:����'��ǟ��S5,���sTM'�61�-D���q��Rcop��kQ�
FwzT0=!�v:'y{$����Դ��w�=��V��ơE�����^����_��U�c�*e�m	-ά��D����m�TI�cO�����n�	ܿ|�ǂ�b��q��s���l�ڴ�Z��q_��EH�.O&����v���w�4��7Z
f��D�l�#/���}N�ٮ�U�:����=9���-H� ��V&��_L�l74�����d;� ן�+\�5�9�]�¢��\�b��F�\�-U�1w�	��aDlʚ[��Ƿ|d*��i�����V�8��\'���y39~�@#�'fz�a��@� �aH��J��M���7��M2{���-\��70�����=������,�3I��nR7�I,�,zn|
�Pe�����/��:��ͧ{�VzI[Qwn�jG�Ʌ ����J]�"]��T���I��7�+<��(1D��\�D+�NG4�L�%^�o0U:�����P�������E���3�otB���@�9� �B(��жD?U��õ��`�gD��o#�d����0v\21����s�d3�����X+�QI;k8Bޜ&����ǳ����e��y�����Ƙ���vXl����E9���6�����va��7�=��2�Bv��Tߺ���/k��\(�����%�6)�u&���{{cv޿�P��x�o�_�(I��r��??Pz�[Nse��a���^��7��3|N�<� �g���!Iey�j��w�B�'Bb����ph��+�Nx@2�����,T����f`�����â�\��|8��JKi��n5qä���i���UT�CEa��4�]"lP��K��V��&S���r�����AY���7��I���	�1��)�|
K�����3�an�>��2��h�3���#�'!^��U���ij(��E��;�Laz�"ӳ��BQ�]���A�)5�L�s��T�Ls1	����m�%˘�N#����g����4~���(+8_t�V�\:uL�|2>�=�3��	ix��K���qm̔آK��;8)r��3�ͽ�M�~�\�'xF�̤E��A�+7�L��kU��sʠ�V�ߎ���{ul_,�]q 7�\�E�hZ�T^f߮���ʩ&��E�^�,�ߴ���S�f�ה�������>$�n���qgS�l�-��g����N|�}Șk߶�V�DsE�����*Ԫ���?2/�;��K��U��\jy��'U3��/o�o������:�&��R�\�RK���Mö�k�8�v����H�� ?T(rf����wiwU���[�TF�И&�9U����	*�����d�Qg�DXP���h�����DC͚���:te����3�ߓ���:v���󫮮�l�ט���:ԕ��u���8-�qӦ��@�4].��f|NĦ�*s8��Iz����:F��xDԔ�6���hb�$��5�9�P��b<e.�@��E�[uf4�*0
���s���i�(d|�w)�M�dwM2���W@)���?�#�e�ܭ��[�)6j���ޑ��a�rc��O�[uf������K�D޲ �e�}�ũwʫY�����!w.��teb�_mX�� Mb���W4�5�9"��֝gl]iۑ� ���A�)�^>G��Z��T6`� �zz���k��xv���Y�(�I<��d�fd�P6P�Qk�2/�y7%����:�:]��Q���ȹ��R_Q>�z�Ӱ�N�~�wJ��s�ߍwDT�6h[\���I��ҹɎ�r���m�ŖE���v���;�T)�X]S�]���vc����#6Jr��dȼ`u���G�j�gq�	�s�|�C���.ՓB��NS�EYt�IQ��!���K����q�(��W�s���I����7�j�7����������t���	�^���7��Ê��}�pG���)�X,w�$�����r�^Lt�pd��\�����ƙ��9$����̩�+�U����j�UD�x�0d��XU��g8Ը�0�����[ID�PL;�_G�#E��sS�bь�A����X����Sv� ]�����v~����wV1ErHk^���n����đyCMowJ7ݠdr�I���Y��§��Fwg�W$�jU�=��dJ��{C�4���}NQ�'�����i��ɚ�}�7����A�3K3p���e�L��c�_��z�0��UDG�ot�R�+q�f��$�~�T�����^0֒��g�A����rs�m��߱��w�����3{�
,n����P�"��L�l����>��t
qW���w�,Q��K"���Esi�h0�	EKE��p���韓��z
T��7��g�ly&Ip0v�_��Z�Q�jqn�7/± �9;����܆�O�[��K��&RHA%�wy�1���l�}�O0k_��'΋-���uE(��T����H3h�|�1#���ct�|˹N=&xփ\R4(�=��1�1@�())�P�gn���մY��0²��cPl�Fz�Q�v��}�fp���3�jȷ�+���7��l��f:N>ʭ�-#�HK٨[����?��a �WO�U�^���-~��w4	,[��&�>� .�P
㩅���L�����嶫T�T0��*K e}V[���"a�5;KjP��d FW���㒊����ʊ�Y�}� {�㻼$��(n�lw���%��C��c�ؠ\��p�h[^I욹HA�����R@�G���3��Ӏ�$�����okdP_x������ۊ�	�uF����ϩH��X�(���3.��sUvQvxq5K ?1Q�+�{I*����Gs���ec1��74���.�������^�MB��A��1�G���RI���ސ�َ݂�J$a�ݸ}C��~iT�͙��u_�Aش�hʆ��>XpndxRu2}��0�Z:��y�����L���Bx����z��*������#Ώ�F� fB��N����_����R�S[��J�DP�+�C�|c�!}wBz�']�zPV~_���K�:�AeX����*��}���?�+OIQ��=p*��
���Ƃ�f�B;P�k�����ϝ�����Ef�~e!��e���7
�������:���I���=*?5��ͻ��t'�#4���B
�go�l�>/*	G;���,y*�����ցf�7�[�� ��j=J�%V�b�=��ѧ�J�v3��1�7܀37H�Y���ɱ|���**8%%e���|9�[3PBd�spi�N������p�|@^cb���4&�36����Ow��磑V�&��4_T�L-���w��|u��&��~�h��^���UZz@�~'\,Ze�7/�^: �"!w���ja��ĲE��'^�����Ra�h��d�qʫ�1=�S��B*;9w&>����-�7�x������=xAv�l�3�_�א��:ǻ��X[��P�%LYǃ������r��Ie�������=��VlA��2���K����Q�M7����0�DWg��<��Qc��S�!�Y�߲��I�Y2���h+g�6�����E"���}�|Co]���"\l���l�5�����*�8A��gM�1����2G���_M�lp/�_�F��`�;�uU���~3�V%?��� ��dJ��6���c�N��n�ڜǣP�>��_��CD�n��-e^�tʹɠ�h���dĝ��גܖ>�#W��6����M�����FQ���_�ꮕ�M
�?|���� ����T�u��=s���|`�چ��V��v�������3�p2��W���V�$�Uy�E{�����l:�<��*Ɛ���(�A.~��WB��A�5j}ghY�~�1.���+�T_L��Z�l�O��خ�<��|�*BW݉�ο6e�8+-	R9pXy=�0��:������b�.[�OJ�脤zc��6����G���qB]�UNf�o��M���Ԑ�;6M������y!����$Ѝ�`�)%��5�a�?�:t���1�ѣ�I�q�#3�?�H�j�Ϫ����j�9���������ysq�5����aD\$��#��ɕh�V�.t�'�Y~�;R���S����c��T�r�P��{]s��������٧>"�?��|��v�ˡU+���n�Cԕ''���8ɁS�3A '�����d�c�P�A�s*���sm4U�V��K#��N������%w��:)L0F�oа4���F�Z��
P���L�U�M��s��ѓ#�O(�g26�6]&N0��I��5���?�!��6'?�nQ-�:,D���+��L_�X��VS��_���C�5E �؅B
��6�a�	�M7�McY7ak�Y�P���X�mˉ��K���%2vë��Нxi�0ߠ�|*_��(W�b�nm֦T�)�7�_Z��W"���x�D߁�,{=�H��?W|V�e��.'�=��y������YtuM\���/��r��Z�E�!�у��>�h�[�5��j3o�:ڋR�O"�l�uoZ���7��g&�rq¸!��|������Y�m����z��������omN7{Sk�r/�*T�r~�*+�J��?�~CW��������P�ʲo�Jw6�ɡԭGrzU�OH���/�M�h8����wL^�������V�^W��=�i�Q�g�q�7����h�՘EI���_��FN�L�^v}�J� ��%t ��a�aY�%-򦶬~��d4C�����x��5o��2Mϛ��Gf|V�M��������+�Z}|�}�����h���>��@��^�C���j���H/a�����<�#��S����m"S�)L�T��3�2O���A��;����rUUmЇ�*�F�/&�P��)TU��<n+:,���>�����Hj�1l��*>p�ĄD��ۚl=�q��2��K�-�y�E0���R�i�Hg ��>՞b�Y�ﶫ���iv��՝��\ѿ΄�Za��,#l >tt�g�̓�zXm�^����f�O����`O��z��A�R_o*�")Q��K��_VD`7�wO�����⎴��j����r�7|�Te��Ff�$�{�7E�X��s��I��ZuKҿ���Ę�.vb��T����:s���#W5[��ݔe�g�81�s������K�K�_�\�%$/jH�O��nΙf.��v�U+�N�����k_�,�]������U�k��/�c|VS|V}}��.�{v�rn�蚬zJ�f��5��԰��";�_	Z�>�H���n�b�<�;|*NӲ��1���@��L�RA�e�a���EjY6V	V�/:�G��*�"g�N���[�W����od��7�:���MI^`q��ԗo@��։M�5
km����2��0P̺
@�IZ0̶���>��l5A�U6����f�<g�8��t����M3s��ZԢ��6%ډ���ʜ���ֶf�����h-ee��/1���_K�vF�8�g����qڝY�p'�zWI5@� zR��eM�K>�T��P��t\��n�sz����%ܿ6����c���i���fO��q�������Ykn<I��@]��m���O�5u��A��Nrb�9��o�e�\t�Zm�x��u��Q!P��][bӃ��ٽ�\��2C��K��J�2;�./�	�f��+�,/[e�,[u���5k?�
��s�}6v$�|*�q��8��^jz�:��=��2���s���k���~�e_���yp�ҷ:��|�tb>�q'@?�NPp��-������T��h�	�g��K���y^P�D2F�}@p-�jOK��Fv������e��g�-]\U`��F��D8�<�1���z��v���u�̢hw^��M�B���:�i��y�-~/,B� ����L��Xޣ�~oc&:����q�s?ێ�q�h�8[ad�"�Cp
D#��x���d�H9�ʮ{�>W2�5���i���^��|
�/�
ְ8=��Kt�v�:rd߆O0|������W�:��#�AC� �tqG׿Q��g-"'[�����긵o�)����:y��S������ ��ܯ��������兼2��m�u�&B��D�$փ2F����!N&�qA����#�K�G����?V�j:���
�:��I�w�����Ȭ�b]0��>��M��??�̥����1��������R���c0ు���m�?����M8�8�ghlE�_�Ə�� AO��z��h�A���O���S�l�H�\��r���4�Cj�B�8�N�с�d\i��4��駔��&�RPo/e��t�XJH��Z,.��8�ԸË���SD7$v�L���X~&�8[N���s̛�#��s��p"�����8���<�FDD��Aj����g˼�saJ[_>�\8�Dj�Ճ�?~������������J$
���NV��w�?���*�(�äƛ7��;(p�?�'����]��W��]�4����U�p�Pp���^�^����ܿt����m]].�C��H�Qؚ��S�;���FH��.!�cpP�Р|)���t�
�gg�$]��K�Ŏ@�H�s@qʡ8�`	YW����5D���۝��ѕ��Α����B��N��O%��N.�445Uon�Ʋ�Щ�$4�������ǅv_��+.C�T�zA)6<��uu�5�ޢ��fU�]$��􋋋ٰ?SCH�� �+��P�/��W�9`��LS~!]���	P"p����k��-#=D�nz��ťW��5��� \܄�.�@6I�1��Z}�����Hc�2{2�WZW3��& � 1P	1J|�j�C�u[�;��@����]3�}��@��M`��o��ӝ�3M�D�C0�Ll��B�|����a��e3`��P�+�d�I��F�9����Sky�h�_�VG�J�b@�6���P|�0�Q9|�:a��]xZ�@H���}�7H���cmm�,BY=1�}o�9��ty�H$�;w���{+dI�Gi��m]������5��+���p^H��e��2b��쬬?DIm��-�t�=,j�f�J`6Ε�iݓ��b���\m����)+�����G�¿a�x��/��vBӄ�B��TPXHOj�V��=��ÇH)6���M����+ߺ�{��Sg�X*2��c:���jj��K�yS��Ǐ��_�jY���j1l�B4��n��ul�^�����4:������G
����}а��|�m�+?�]�?0���XtJ���3R���+��Gܿ)�hhj�K��(��3�3m�=@0i�jbb�+�A�O=Gy`�
�!��Qb\|�bG������O�<����
I�3}��
�"w�<�G�m�:l��>^��T��펙�|���&W��ɾXۏA[2��h4��RM�3^��\b�M�W��8�}����	��[�����<�Y/)$o0	��p�S�2�pLj(@F��$�l��Ҧ:v,���6��klj
��ӛoc����q�%C����BA�*���~On]x��YZ�~�f��i{���^�vs� ���h�&T�0�����w�=|��C�Q�iM�W��?2}�O2W�X^�G���������R?@�W�Y~5���Zd�PAMԑ���9�}?�h-�}cEk`������BC\{�Y���֩n]�A� ujr��Y�,oƴy�aIMZ�k
�Tq,{�P�	�+~+нl���l�(�����l�9��I��|$�w�@r9��m�_'�ꨧ3YW��<J���+����=]�}}��F���~�����a��	�\8z&&�ngN�N�)P3힚-���*�����ع����8�-�F-�빜Ej��6w�nі%�.
q^ӽ��������:����T �8f	�
[n�+���(���d<��m���K�����-�{X3f�82����T�[W��\�|��5�t��3�6���D5�_Yzz�������h�*�-5�8Ja��t%))I��Iz�W��o�ځ��{����S`d�>N�(U+M.��~|��U��Dr75y�P��!w�=G3�>6��Dl����}�cg$ �o;Ȭ�o}9[U�ƍ�-�#-��$�Mhp��:4�e{�	:7��'�(?��܄��%�E͊ڏ?��2�p�բ�<�9ML����F��^6��c"}|���RS^ZX�j��~A�b���J#F���l�qUS�O�mll4p~����� ua͕��s7��m���%����q�HY���3�ֿt瘛8����+X�>U��E״����g�j�A[��]䞣�[����y��`��V��H�C�i��A��#,F���z��W�,J�F�����Ề��:k��7n�8WfY�]�6}e{444t�������ޮ�q�aS�� �N/��.����ȷ�n��6��{l���3R�x�,h��u�P�Y����4��M�g��w���˿+��q��G"�^I����٘��c�^�)��f���A���P�R�hS�8��Ӈ�
�|1�ف�����1i�ò	6���=�Q��{�p�&���T���� +���F���l�L[��q��=w�v����ʰ֘�^^>�j8�=sʚ楯�oW�����~��`7���P���p.j�IF�(�<�z:�f��?TU�2^��K'+��<���e��Aq�����ZXI����{�(�~��_M���o��q�t�W"R�д�G��r���P�.)}� O���j	8��gce�WP0�X]Sc��\D�uez�&DI���fH�F��ٗQQ�e��|׆�Qt��?�c��8P���C�jum�H_6;7׾�H�ҥ���rM��R��!8���W��H��(�����ӞNߎU��)��*����O�	dڨϧ98n�G�Ke�`��1����� |X�F�yHH@�Vm$y����9pBd�o�)(!���s�y�x4��zxH�ٞ�C�)����"�	l헮W�����8͕X�i��c�U�%���(��h�9=��]������	�y*�6S�|d&�����A��A.���WD���?)�}�?��\'*����=�:�-wnR��ǟ�J����$>�= �v`���A@�+�)b��X䈷�wɫ��
7//�G�<||��zy����if���x��M�%,I3�b%����ͬE>Y%���Z��/(C��pۚ2
J�q�BWl�n��&�:�>a�Ɍe�i��9�}���� �r@���
����gzŁ��LR�VV�|��:LWA�*�v/�j0�+���Nc����8�o���r�S����qP�ִ��e�"��և~}�p�ɩ0�$�)�� V%�*)�
�+b�DV�HRt��	�g
��&�؁|$� .�E<��
pi�(�D3O7���..&�N6�X��<m�z^��׍vUi&�U��Sˬ���AQ���r���l�`��Fڗ@�O�
��,g���l2����
��9�*�j�IM`W�+�w#+���{��L43U��w7*�%��V�dYq���� 0���Y���p�豞�)�i11q#H��3���[W�2ɓxPR��s����S�{j�n��j�Ν����1W���	�q�	b�п{E��{�;�i�$���t3��[��Fku�Ť
N��H���٨`�uܸko���>�9E�)���A&�I,-�`
�z���r�>(��2�Eث
����rF�XܗZcx2E�cʛ_Y�� �6��5U�QZ΢�
����Z�,�:��p���i�p�:��$�W�����H�u�LYm/��1�4��+fH��6QP ���2�\[��hXP:ʛr��[f�&i�-�����*��Gq��.i�B���(Y��O-6K�x��{v�F���j
��]��g�Μy����4�7xFd���?((<о��z�ʝ�Ov�8=2����Y<�s��q��@�4s2��6~�+0;�Ñ��}JO�"��:��@a϶�5���er�.+�qG����\����é
\�������"��G4R�t��ߺJU\��Q����";'�7��]!		Ɛ��#"�7D�O �O�c6n3T��b�kmW�þ����ʩ�X��n��nsq��A����{Dr�YUa, (H!Ow�>`u�^����w�d(wA� G�{��;�Z[[i�͒ѮI4�^=+��Z+-�{`�.�;o�B��+�azh_�h6��jO�CQ77�z���_(4�ū��;7g����� �T�t8e�<H�]@��q�Cũ�����fgg6�/J�,jkk�w��1��ǯQJӃ�4�D>�7��eh���%b��o�h�RK���t����"[��E�VZf�R��CUu��c:S���ty�]�e6L�U��R�jM��`ߊ��ȈM��/4�Ȗy��V�W���%|	�e�)+�	F�L���E��E1M����Sy��l9ŵ�+ֿ8��8�b�%`���O��4E����^��������0���� ��:���͕(�U�^�ZO�.eRv���p���T8��#eU�r�aאpK�\a�3x�S���,�)�;4���$�:�ye�����i�#���߹����HQv�u[���~�����=�<|\��g�c�E�P��,���R$�4g��V.l���1����G��F��{�O� >J'}��W A8<�L�z6�Zr#�Y]�_��s-�4׿���������֜�?��J%G���{P��E[ME (�Z�G�Ib��c�^ށ}�,
К���ͷ�B��\�Ə�r� �fcc���oS���ވB����eC��� ���*��4Ѫ��+ߵ�Le#;lq�6P��48�HhӁ��i� �cy������Cp���h:���7�(W��?J �1�;V��Yafd��(jQ:�e��x[N@�,�k?����s5ˍ�pC��i!�w  �Y��tog�(�I���>lS���&����l��
����V����2K{����C
�_�x�m�4777����<q��ի�S}���Ĩ=�O��:�)Ж^�>�_&��)6�RSTV��-9O��y�}���|)��h'��4;�w�@�v�[3&�&&q��8��Lh�u1��-��-����n5)4��𭷀+=�/�*
N�j���:�Jԕ�L�#����5�B�_���n���N%����Eח��th�o���YҦ5AmM5�d�\�{B�E�kK��90�9��B'�&���#u���ᗫ��Wb�j���B�Cň��R�C��SU�w�.�'�d��M��TWWGv&3���f1M��$%�,.�QPQ���#3��^�Z�����R2^W$���o�|AEIa¬�v>VEC�b1��q^]�Y$\;p����Oh]9]��m����6��f׸����e��8&u|��H�9ݛ���y'7�#UF1��Zb�P?���a�����=w�Azjs]�J�ͪ}�n��e�%:ZQV-����:ʜ�cQ$�a�]7٨f�X����!�ta�Gh��lfJ���;�cVf�{�.��
򱕯:N;�ִ��ǉ�`���Դ�J�AL�u�̄nkC2i��Hh�[w{��H� ��D<s���n�s���չ���w�ٿ�s�\F�ž|�`�@�q}4*6��k/̀ei#����!�K�0��`�h�v$%$6�>x���0�e�#˽nRB��^Ʒ��ȐI�"�i�8��@:w�e����\z�<ϻM�#�v�`��+�����ߡ\�s%�J�VT|^��Y���\YZZ�V����XU�\�qD��ɌW(5�Su�y��	��BC��|p��[>VC�x����N��:���:1QzH����Cޑ�bA)���ߗ�m���d�qN��#�:h�����=yi�#� *,b�qo�]�B���n�S���'�Ѕ������|J؆)C{�_Ft��� �8��ɺٹ��?w�9腾�a��`�%�Ӗ��o�Ҥ_�QW�ENW^��b�gPC�)t �i�~�H����x�X0rmm�#S��W�,�VP���@���S�"�,i�� �X��K�Q��8�n܈<�_G�.��l{��V��J�I���Ev����
��;m�o�x_)�\��B�e��_���3b���נ�Os4��?;{J_�r�!��N�7�_�X����j�D��;�T�rF3+#��*u�CHfj����eي0���y'�>j(��3���g(ՔG�x.����*QRTʑ�s����"�a��H���Z�(�-�G���lT��Z�wq-�U<�%���b�����/i�\ G��`�����>z7D�t�`%�E����w��O�}}�c@�j�?�ܗ��{�i�|g�'�UG�dRKT�{�+B̏�өl�B<��6����9��y������sǊ �k=�@�5�2C���b�d�����rٗ��)����S�퀌=�>NN���7�d0����/aAĝꩩ�rgL��(pg�;��%ќz}J7A����o��V�y+s�`��[��B���������Z��Q�J3�Y� KY���3_f�E~_k�N�uԄ��^�$�n�(��V1��8�� ,�2��bp�������w�y@��+J(�9�T2�gjb��ȩ�嚯���@�%z*V�}�H�q��C�HSP())�7�N�d8�
��}�@�b�T���P\(wgY'����Z}Lg����;���w|_�+������C�6;?�q�?j���P�q��[T�	���&Ȃ�Z][�<�U�C���;&��^a<uVP A�q� �u�;&��B���m�X!5ԹW���E�1��~�HGg��Gw	VL��~��Z���|^^�$�s�Wy�����`�)��e�^k�C��H�B@:�|G B�\���l��q:@�uj%�w�w�--e�3�:�\�1%�w�w��tO�2V�b�Nþ�'�b� -�g��x5�"�9`����*�z���tck��a��۲EZ����H�\~A�	�ls������L�� ��GHx���]RXDď4ekck[Q�x�laZ8::�h~)q��b�@��H=��� x&�,8�����1���$E<I;��S3MK����:5݌9��Z<���鮾����,.˓�<,�W>T�ih��7
	��V�s�_V6f�j�BxhCz�n�bj���h]���KNƒ���Fl���i[pmJ��p~M͜�EU==�
�)(�a��g 8�Z����"��EG-
���d�֘��N�
p�윜��ME�C�/F���2S����+���)��yצū�7�|����uH5�-��KIm�-��!�]����za}k��<��V1�S;��6��r��Ba|�.e���o߶U-fv8l�4K��</�_�P�) ����]���#d��hJJJ�H.hN+��ut|�uu-�V�E-��82u#l���jzzt�5<���M�Q��Y,��7l�or��XR����cu��ϊ��P�{�
 'LĿ�8A���VZ0By�t�j1����y��������ԗ؞h�'��{Z�B�O�W����"�ʥ��8:9��&�A�t'ڦ�_�VZT@;�&�O�S����q+q��3��Y&h�Bu�u��08`s�k=��e�^�ٿf$�r�!hU�7o����TVAlZ��⌄�	ق� ���jRqFd��)Q֘���������׬�uR��dJ�/X�"3�QI�Cn�6t"m
�H���� $��q�S�אs�R:�_hNPT�a��Q/9GV�)P��J����/����8�ֈ}�:iNCM�6�r�JM�{sT��m�v~~���	�):�}'�}VRS=F���F��A�$�Du)��HSs�8��� ���[�z������&�/��10gN. c�]�����1?"�)3K�(U^�Q@x$^K]%	K�KjF���H�8y��@���ylՙя�pE�CȎ�O�l��T#Yt!d�d�~|�7��4�R?:#�y��ǐ�,v���X�aY�Yǒخ�ޒ^{N(�1L�w/'�"�g�������"���o����I����ooo#����B'F� ~�UgQ���	{�"���,���vG�]���%�&f����RX�d7e�%/���i�Gδ
�O,���Ǩ�H�����>��6�V�a0�)P��L�˿X� .vgx�u�6ۜܟ���l�����?PK   |G�X�v��f �� /   images/153184b0-233d-45e0-a203-5756afb39f29.jpg�|w U�������JF7��\;�F$�Uff�����M������$���k�l23�M��{�T�|����߹����>��<����sn�} ͅ�
�  ���
�����������|QS�`T�h�������������	s�8�),!�/(�x����{<���e�>R"� ���}�}���� � � ���FH% ������ PB"�N F �hh  ��M.`�����l|�W�	����w���g ����v�9��Y?m$W�WV3�2�K��5�Wh�F��x����v�FI�d��UaV�k��Z��o�����
��s�g�ǆ���18��61QG6s�E̖��x�*�ގ���Rymd�2��S�zj������-S]t�8��֚:b�.�:Z���
�ޛ�]GdT��4$�I(�N�b��C�y6 �^��r�>z�W>�L;T9��u�,���&���XarEU��o��jwj��"�.y�B5�cjɩ��Cfe~�~q#�y]���e�7M9S6_Um`�\M�,_��%�ܓ��k3O��|�[�}�����K|Wf������ ��smS����~�����bw,�3{��#�I�\�m�{�SK�ĵqn���ś��j����[��Y��|�nQ�5m�q��՝�J�q�$W㞉S�<g��>.��=�A�ϣ�Ԯ��PGc�qq���bW�V��-�6=l���b#�[ b�
�;f��şx�������T����B�-k�56�#-�aK���uS�>f���w���׌�;O6�l~%�����/�Y��P��L ���k(�mx��\ �f�ጥ:F"6 Xr|�P���3���X����	�47[[*�n�J��J5�]���1�Ųo��d�wbz�#kK�Zf]��R����^z-��򴹽M{�q:hB��xe�B��t�!ͻ������n�$�[��NF����YC�����~�1f-��w���Z�+����/�5F�.*I���~~ڝ�Ʊ7��K�� S�k�c�1����Q��.$�-�@G�c�y�nx��9�Nr��D�O��D�U��x'�(���Ŷ^��B���!'-�cɝ��>��)PՅx-�
������".N��
��t�[=	O�V�?)r�!{���`�mG�`R���۰Յ=s�i��z��zw4��b�|�]�����f�0��9� ��Q��KY�7y����e%"��L�x��R��Dv�����>�۲Іy��٘"F=Qm�Qш{�L�[Ɏ�N6���KC�nW�0�/�/|��M!+iL*C[���<��g�I��ZB���Ʈ�]���ۭo��\��_ܙI:Q��T��)�;V)<r_���G#���B}2��Y9�9֚Ƶǻu���M���=�r��9��'��Kl�>�E���兄�h|��M���?�F�������J�gϟ�������/]s��D>1QS�����)��;�����G�mX��CI�o�Qˠx�?����;�����Y��G��JW���rZx'Tj�pc�H7&�`q�X�X
\�Ngy�MR�*����|��0m�	����o8FU=�6r7���5;��*����1��:w��ۀY�3��
C��#����}��K��� Z!�lЭm��"}?}r]�h9i���97��r�k��H��=�Rt\���� I�ʸ��5W��Ob�=(2d�Z�`�_���DF�8 ��PG�l�;��x��?� �}�z��x��6�^&�%�r���qA��KEk�������/��9���髃���O�6v*�
�:�?	�%�K���縹���J��[���3m f��93��{�)�zי��y���{��BW�`eR&<��B�X��3M����x�x�7�S�e_��.�w�����_��p΋B�D��۞��FJ��N�W�/:\�w?;5��N�T�|Dg�,����Q�r��b�{@��ǳ�������ht:/cafV��~>�={) �>��Dн�{�9:��|e2���B{hpF�.9�-��)x<]B<eKb���	��a{���"K�-pgڇ��';����M|(9�Uy��Q�m�8p��,��%���-�`�z��G��C{�w�)a��3w�d���h���~S�8g���F*�N=�f�"#���q��s���hD���t��N�F�>�㣌?R�N��Z6�� ���������#�>�ҷ8�uj-ݝ�sn�)�Ze�/���_v�����l#�Hi䜮wp�"�<���}kyؘhI��HU�K%h���Pp�9���(�����|�j�s.&�,�sןǲ��4K���b�t�#Z��|-�}|*$Eu-�'v4����m�y��h��:��E�k�Ln���u�y�p��Z�@P���J��z�i�3���A�[�u~��S�w��<pazsk�'>ky�j�K�ܟ%�x�x���������Bh�4�������k�o��~��f�t3��fO���c���hB���������K�?H.>_;��>I�7�hv���I�n��ec�ޒ�v����~X��C���w�y��1��Q(����8�n��P�j�pn	�[3����Y7�{q�@�D�"�{f2�Aj+�%�[Y\���Mf�V�>�m�
Ӯd.�,��8�b�=(��,.�'�$h{{m��3Ih�a9)�W%_�g�g�lk([�)��������ݴ*�h��+7;�<����9��.l�Ѡ}[t�,�e���u~ݓpș��[����y�ٳ~ұA�z��-���&�k�����	t�T�.Yn��Ng����}��O���Q쨭���W�+R9C���.���R�͢*�K����L�UY�<;��gI�#�w>[�h�E�F+=h����B�;��������[8�ώᶈc�x��&�Y�Q�ڏ!4�th.�IďǏ#� ��-<m��9�XW릢�_������=�/�|12�|�{�O|=�$�8~X45�'=�Q���vo� �4�Ϛ�l(��:�٠�C�A����Y3�H��9?	�.�<��n���P.�妗�� �}lr�R[߇ՅSw_�a���*c�1^f|���:�����X\g�wrK�����J��{ȱ��U�3&
��ܣ��\L}M�R�^�d �Փu?�ĩ+4I~{�4���F��s�����LbU$��Gn�ЅX�d�"��ʛ_s�;���N9^qmIe��f
�"�u;ʽn]��?�1� 
�=Þ�v'� ��wѡ>!�2��}w�)�Y�L��g�g�(��=+A��ؾ"TO�,22�o�Ag+��x�=]�Sh���������V*��p��u!��2^�<���pQ
�ϥ�~vY��_�T����|g�9mi��zS�Z9�wk3�}�M�/vjى�;>Rxn�Y�A�ˍ�:��`O�R��=+m���f&>ԝ�ݚ�/%��̗��`�����Оo���Vφ���wr8��;�H�ųw��-���*��qQ��"8q�����\#��pǾ�Zv����Z�2�ωt5�	�.��q������G�0��dj8Ы�{�Vd}E�:Ύ��%�~.<�赩]y�t���#�����ca'5I$��nE��+&ԒN�u>�OE���H�&_+�|w��P��Z��_py'��x>P�gP�����m^�e��Re��0����[��{\V�P.�3iA�g���7G�#O;*<;���ϭE���CK.�M����^,�3ċF�&Xr�[<6%n�ì����Lp�T{B^RN��������Ю�'�C�*?�{�W�c�<�1�[4�5z��T���T���v�w�9!�Q;E��{��$���q�� �4���!Q���y����
Z��CGl�p�n�](@��"���O�zS}Ƶ1[������mp] >�6`�b��Ȏ�y�g���^gI1���Ù�`�H�ÒK�.���j�I*�V�eJώ�9�Q�\� ���3����3�_&1q��M����� ��wz 	#w{���p����n�������ȩ|f����U�#�ΰ�����'���1zڨ5lg��M�9M���dH�"{�^�ڵ�VEvP=ͥDU��3�����u�fSݚo\��;�+�����vGQ�*.5�ՙ�5��j�m��?�H���/�v�6+N�� _M���DH�b��QE�O`�Jl�.���^��m�u��ë��++�W�������;uF3��!�G���ddZ��(wolðh������{��;8�0-g�AL�ǵ^�Uz�N���El�������#�RPv:9�2dĿ��]嵴H��b��!#h����c~���-�T��Y`�u�������-�{'������7�����2�2��DF�X���T�����t��w��"n��y6��b{��m^^ �n\s���52��#��gN>�[7δ�9��3.�M3���͛'�4�~ߓ�.�Su>(��^���x�Ģú�Y�"�l�7��W�.�AGVqt����\�qsڐ�*\�j#^*T*�3V�}ߌ�=O�V�Ix�ȵ0��;f�$[�u�GD�).ݤ�I0�k}Se�l���2�}Ҭ���4�!�^� V�ZP���f-��c�1�&1)J��$�Q���Fȥ����t���Iϲ�3x�ՏMǎ���Nގ���:8�|�F�>N�MZ��s���[SK�z��'�Jb#��1-9�/�`�;�X% ��(�$P�m�0�u�Z`^W�����'r��OO^���9�!����Y�ף�b�<�\2����������.���R����+3ײ2�����
#p�sSG�RX?��E�*��S+ �x��!h�g�����d�j�'��(� K�#W���>� ���x̽�c|;���'�z�)��r.5�"��^7��Ƭ�ާ8�Z�'2(�M��`�XN��ࠡ����n]#������\�!���:غq���
\�S��������s�*ʐ=f�Y��PJ��õZt��(�4�`K�ɍ�v�³iT͇�KÓ�<S#���K7�U�����w{�8'���/�������\��t�h��X����~�~Qͺ��ت�[H�k�'#��Z�0��*4tZ<<!q�B�ira�%���=�'cfn2u
�ȧ&(��GҏOj���k`G�]a�}�WWz�����/����y�Yh�nO�X���+r^]�q��ud{�h�^|����0Tk{�fi4��D�ِh
��bˎu�K'[�k�q�ŗF ���u�˴xt��؍���ĩ=�[]Wl;'����Ɓy�wIZoZ�҅��[m 烖n���3�H����휔���^*��1�Q1�v�lqq
�-�	Ig5��q�}P�# �k#2�m����Vy��O�.�ߩ��/��	p�8x|;6o���V՞?ݗ�n�``f���J�i�c��r,�;�]/K�7��%͎����9B��ߛ���'���-��<Ṩ-`yH��Q�F�)P$�C�_���KX/�r��jHMQl�y��݂�u>A��(T�r=j�0�{�](�.�QV��DG����,�y'�����>�п��]��
Oy5h@����~x2��͝�'�JO��Ta~���c�l��ʼ~t�-��\G�C�vo�K�T7gZD�j����M�Ґ�2��7����4N	��aG��IʟmM/>�n�j��q ������wX� c��L�����J�=]���o��|����3'���d�z���QL�+,��M���t��U�j�Ic����B��H��2�f^� #�	I]�X~DzH�s.����<0�,��U�n��XG6]�\%�5�8�2'�֬�F �k>,ob�)"uT�����"��;R �S=e��kf~�5R����h��%�GɪfZ���� O�1�e)��S�����it��n����Hu�|v�k��l��Xӛ�_]�v05CS�vqtam���=�a9���v�%�y��z�qM1_��~��� ��;b&��}������dT��#���àoyB�=�7�=ᣀ��'� ��qr���)W|]z8F���e����j#��ް��Nn߂�Uj��#��p�;��ON��p=nܫ�&�w����W�.�W�}��E��&f�b]���_g�ԫ�@��=�o&|���'��B����"��e���6���cJnd�J���I�/��y��&�?j�����;��.)���AF�!�	S�
%_�������u��91�↶��Q�]*�� \ �*�@c���;�+m���gN�G������
\� a��~��P��%���.9�}��%E���W�b�|�,m?#�S �.\vma]$x΅d�'r(/�����[r؂,�w������}��H�:��3b�	AF���j+>��T�o�v�$�.�D�B�}rX�ĥ7�S�n����9�t:_
�D�ΠÂ1Tg�\��'3��!$O�|��	���f�����I��Iy����w� �h�������!�rM3����|�K���w��Õ���V|�	�2-��G�_�a^��������V��Pw�;\�l�g�ǷbyԜ�p�o��V�u��������y�!���� �R+��ೕK��˳�sf�ܿn�'�;=��+|0�vX��LtD����e_g�m�z�%-$�k:b�� ;hb%�K�偉�ۀ��Q�j����uj,&�����LA�J�'q;"����E�F�PKa.�-��֓��y�={4ۑ��t�F��W0�[�B�/|X-b�V��{F�Q��J���fn3����_�*>�+^��axC\���}����CRl��"��Fc��䄎��JȮ����b/~]8���eNo�n}����Б�́�Tst	��[�3����.��,ޒ�2����h���f�>���AV�6����`�Z�'-GSl�,+�Qw�҆ץ�����k�?�R��&���Z��8�g��h�8��5��,����r;��cg�M�4#-u;����o���G�� ���� �;RlB�}��v{,��@���8w��S�l�d�[���f��.���F|��VP�>�qy{��E��^�-����,�N��n��L�5p>aw�)��4���9��$���,^6��O�E�N�I���_cjJ�F��G��(��C�w�a;�[c`?�h����`S��3ǹJ�x�����THw��z˒�7{�=��%�.���Y�q�mz�3�B!��g��U廒�u��ϊ���}��en��[�U�����]�;D9�;Gb�n6w
	?�냟���sc�n̏�O�i�f�p��]��Z^f�Pp?W�ؾ�{7�y������rl�_���,�it^2�[�ޝ�4ߚ���k ���г �[�T?|����� L��7��_��i!'Cy��l������'ɱ�;��݌6�K���r�4NÕd�-�����@<�u��\��	��54H�p����G���#P�� D�-  ��	�H�]�����!��>��k�nd���htt��3�����:�,|�������q?�V;�Ϙ����~���ʩ!���E���������CdiǊ���;?�\{�\��i�o�"r��U������x�r�]n�Rx6P{����ZåI�{��[Qp���?���֯��N��V��h��L@Y$��B6����@�*õ�-�6]����XL����|�~�� ���3E�v�.�髭53ҋN/:��V��4-�ʏۉ������dsc7v�
��Nz�z�dr1]��N�+���^!���Z�cN^2h�f��m���?�@[�sl�c�%���(��[;�����R�x��~���E(�OGZ�(���P���]��|`�����FvP,��"����Fv��k�X�<���?a2��to���C�Wq��SǄ�H6(ֿ������3�~!���W���z�O5t�%����a���N��v;�1����k�����&;~���\�C�����#(Vٺ���
�TK�����R��̴�^ydm��P��=�ݨ��Ii��DV4l���C(�-�A
��A+?{��q�׽� �f��c�|��m�Y)ӗ�*%7N��^8�qI&x>q`K9��S��M%��M�Ό�j��V��(�0���ۆ�N�1�����(%3�8sR �D����/�"%~>a̱�֒s�k -sv�2G�V��c$�
1���+K=·�9T_��&�\�9����6T~@��ɡC(����ڳY��w�o�D��S��{4���������W�	b�Lm�v�u�ا�O�cW����wp�t?�.�mxn"Oa�U݋Xf��� �*����X���7�^��� k5�!����J��Wf�j�C����F�rhZ��T�:a�`<�L�I�պ���rf���
Sݫ�5hJ�BuЉ|!�_���dnF[[�\��f��rʂo�ώĈ�X��|²Ud��K� ������yծ������1�ة�W"�!��wG��N�;-8N|H�e�(� �L�#�$�+4F`�_���Sj�� �Wƭ�p6�����+e�����O�C�n+\�
��Y�&׽#C�]��%�fWh�%I�?���]�x&��H�p#u��3E<�Tn�+���[9_���V.�.<��#�������2+lp'/Yu�;w[E���cNZ�v��M���T�~
��
�v��	�gu�ƕB���q�#��|��TrS�H�������iΟ;+��7rh>����f�?�����we�<H��ܳ7L^�o�vA7g��v�
oz��~�ȵ˧�ށI��M�dS+��+Z�^O2�ʔ/t�p>!R`"%���/	���K<���Vy�o�<ɦ��䱐����]ï'��8����y[���j*�o,Ň�̩�<�J�����J�
n�ӷ��#�;���0�"�b�f����`��Є����V�#�P�N��[�	��G'�H���� 噜0���-$6�R��+d��%]w9vG(��J ���'�v���V����)W��qQ���9�)�3��5u*�L���hE<��w(
��7�2}2 �qŜw�����si����(�C��V"�ɗ�S��N��U��υ�Z�q���#���T/6\M?p8���fi�/�w�q���g�}D�T�����ؼ���rj[�W�ȗ(a��U@alypNm8���v{ �c��1����讖��U[I��iS��K�x�wަCN�79����[�m�ǔ�_����멺?�a�^�k���X��R;���_hM+߾U��FV}sP
;e{�-�y��V#
h*T@yH����TX��a�*�,��cC��F��_�AgG�Mm~?�X>��n�z3\ ����}ƾ�]�v��#��-�y��6���o{�~�>=J�a<Y9��,�[��y�E��h{߀<I�1p�� ���Bc޽?n��dӐHgO�HՒѬۈ_�8��~��)/"�S�r���Jܽ���y����i��u<�	�,���<"0qB����$*� �F�P�AXc��j, �v���C/ǠbR����Hw>��ݤ*@�1����ue�	����+?_��_�d'X-5�l�ͱ����#c��7j�`��.�W��g���A�x�M���T�Y���#|�M�ߔ�����g�bY�>�����QC���(���~Y��v���z�
��w��g�a��w����ʖa\�\�#�׌���a�i����i�!*'擣/�e�rN�<�l�0Ӓ���R����F�/�b�~����C�UZ�F�kn����*X�Լ�l�"_������w�����_�E
��YԢ���>K<�7_doˋ��]��NRk�O�*h�U Dݕ ����A=����|v�;�PWɠ��ޕюa%3g��.KJN7�3/l^���n�]��"����u_Ԓ�(�W�b������b�0����o�[�fifh7V-�,L{w,P�0J��h��H���H��(K.^���?f�p<��b	�5s/Dͦ�fb�����vO����(j�Fخf�Ӥ���p�$R4/�n��\@-���Q��;g&��7�<'�c���(�K+f��?����`�{�!qƟ���z?�������I) ����6l9�yQ}�|��kaU�����Q@p6�W}�Q��2��Fо�y�o���d�4��n<1����ĩq��w�1Y�g�j�#�ۊ7��!�.�'W�"�A�XL�:v"���������cv�"�
���68p,p �S�F��A�m�
����kC��:HL�𤷒������ �g#�r��2u�G@��᯼/:?.f6�fD|�}���C�M߾��:����n4�֥���n%"L���&�{��;b[�����qJx.�zNPK��X��k\Ö<��	��*�p�N�;z��]��$�{A?t���L(O���H媸=M�ơ X��%�L�\@�!��X�3 9��^;�T�N����[&��E�`=���G��WYq�	��CK{�]�D ,t�r~譳��� ����4b=��.OU�.`�5q�v�,�j1t8lH$�P���H�3]�_*���t����&�{'Ğl�^KK�̀3J��m/$�������ph&�<�G���\�#Ӈ�cd���>�K!AV����K�)�3�����X�]����!���\��#O�24�t�X7�%ɕ���� ��4��,~Z��g�>�3�k���l�#�
��p{����F{����T�]�K������8WA����I� rA�Z;�H��K5�,��i�}�L�4d�=-�:�{G�������@�}y�/�ݻ)����D��|mhq������~&���H��ÿb��l:W8W�[���Т ��]
㖫�8��U������[g��pu��.>u].`X�Ј +�r�F"������a.@;���H{-�@�g�\�φ'%E���m��5�69�<�����]��	�0�B吨D)I$�ާ����LQ�l����|�6k�Y~�DD��k�Y��3I�<�I⥶�A�|�{e3ŢZ�D��l��W-g��J.aFG�;��;ّ�M�L��m3��i*��,�3,���.��+����|E���o�oW�b��Z���+���Ly|��rD�ƚQy��o�cX�E����"3'_�cW��7�<���Ǿ�ӂ�%�:Ipr���X5a���X�{����,�HW�<��x� ��g�6M�r�g]�����?#/�4҃#Ǻa������2�W�)K�̻r��'8� R�Yp�a�\�4ˡ�$p�����2?ҙ�%���͋nR��jL*�BŒ���GY�d�$���T�;�w�# ���!@��Smh�/7)���BĖ���B#��0�ߤq����\�K�yu�՛�ȴ�(:,�Bv�hC���U>�V6I����YL�� �uYP�T��+s-�������)󶤠�~�q����dl��Ԓ,.������
8~��ƭ�P�>�g�@��R�* QcES���5v�!���`��C��4��>e���(�X"�*�h/�*8�}�:E��\�5cx+�H��)
 ��i@��UA� 2  ����A9 ��������֣�j�>��R����wh�i���`H��c:�Ej����*�����8D��[h�7Q�a�Z��(�9����,@����1 N�����6�%�����k�`�Ja4�Pď��� ��{��������d������yRwz�a߿��ӥ�t��X�sB�dB8
�%���;�)���S���!@�	z?�5;��|�(�U�J1�;Ii�	^��[y)loɵ���M^� -�����@v�-X�V
��L\n��p~{N�<�/���#�=v�y Ρؤ�K)����-���W2�\weP_Q�c�[�y���-j�y&0'��[���� �g��(�;$L(M�'v� Υ���!�G� �js�p&���!��
���t02��r ��4�i- g�L�֭�l�_h8�.ݷΒd�5�z���Q�5"U��J��RLm���G1(e�m%�(u�OG�d�[JU@���e�<m� �=� 'Zvt�gqsJ�>KHs�����Y�	�dC���z���'����3�O&��ί�e�~B�/�GFu[<צ��H�Q���kHB��%��U(��p��@l�Ȩ�%�&�ӛJ���)�� �OG��&�!��^u��:�*HD�z9nLf���3�>ƨl�Az� �覗�T�N�S�F��,�qQ��2�m�	w��t�lR�)���9"|4GI_;�%k����.'���+�.5x=��/Hm�[�pgU�F����EH=Ȟ�}ٛ��z7�M�|�� �Tc%8� �>;�Z�5))�pl��}td�r�TS�� �"9�@�ck)�Ώ���Q;�	"ݐ�p8�Ԙ���=?$vq?H=]\O͎�����hPf��jǷ�fd��<�.�J������D9�2�����y��A��r6%7Մ�f����zL"��#H�g%��Mx�%��(?�c���?T�v]�1�@N�,IVX�n��,���&p���?����r:�&t��Q�d�q�dh�Y\l�q����WӀz������o��������}�Q��1V�d2}o��!a2��'mxrGy���ߖʬMo�L̄��=�:K�4��(E�9��Ğ��N �S�CfrR@勪���)
9���,!��:~���`�@39Q:��}���n��6�˷.���D�<�D���=�%�U
�����PI: Q�ܢ�A�u�tj+v����`8օ��������:��-Pn�Mp0
s�G�܀j��d�,U0��l�)�0���c����Y��V�i�`�~�r!28��w�1SC�;h��6�)�y�;��\s��#;�m�g@���9���r�=�Yp:��N?���dT��b:}������h��pP�(H�iSF�2��(�_`\ģ�=�å[[�}��`��"� ��$���(藬�_=#�\�V)SX�R�	��B+lQd�G\���H��b.� �T�� �ޢ�
D�4�Ī?^wL��h��GF)�,�%�p������2� �:]_ �m�7�lfa�̡���_�k�S�R�H�`��L٥������_`�N|��L[�zVye�i�<�W��o5-=��b�tH����k�(Di��啼 ߃xx#���q����c4�x T��� k'Ie|O�^�UD�(��.�+ �����m̥��X�����xD�}"�_P��s�H��5PtEP_nX�k��W2 \����r�.lϛ\�e�Z
���]�5F��6���W*�����Z=�Bs�����6���0��tY!JȨ=��)�&��,�5��gܶ�:]d���X,��&B���{�K�绛���)�h����aNK�?z#���o�=��,���uj�����o�_X����5n�f�:xo���*�c��a뜤�XJ� d/���%�X�4��	�*��s5}��SA��L����5�pn5��/tDV57�sMԽ�ǥ�@.\���c�َ��J�� [iyXg·�gQ X���m�¾���N��� � �Bu���щW�z�w�.�~�)�M�nQG=b�!`Ҥ �^���Q���MڛQ]
@��K��E�"���Yb�;Ӟ=E��K]��zԁ�ƅ ��K��&62�1��rr�4 �ś�+J D%j��ϢD ��{�t,L���Y��7(����]�T�Fm��Ji (wV|��Y6�Wʦ��G����aϐ����|��Kvm4^���0@&*ǃ;B�p�ӄ*���X8��*9� ���
:O�e�d[�?ݵ��}��k�fY���!鵇�W�p;+n���!i����_{T.����SJQ=Q�Hd,!�%�t�M���n�K �ϟ����=|����@���Xm�z�c�wf2�Q����������~��qWB�	��������|x�h���a��J�� ��45U,�-�י:�^)�tG���R��|�z��{#2=��>28R�j��d���Z)u�� �+���ǰ,ͯ��� ��6�o�ȹf�O�i�����p#.~��Rh���w=���]�����p�}v�^���z�('C4�c)j�c�J
w��Sb��[g��D��-�}\�����gy��gQ{`�����;s���`�a�x��<���r��dE�:է��{�`	��(��M���e����@ܮV�^t������%�l�`�+��s�-b�������5�_�ꟑM�^����VC�P�ԋb��rFL�}[_�m��yQ����v���r�k0����3��#��A0X���6�D�4�k_G��˪cj��@,L
�E"Mc\�E���'v��(-E)�ӗ�Т���6V�����>X���7�!;�$g�ڴ�դ+��H���6V�؃)��<N�2 �V�vFI&'T�����{9M	lc0h�qաc�^4�����U��m 
��N��ώ�`I �Z��T_��)Yq����H�dLCh�
J\J�0�ź��0p���g �3V���� D��f%)(2���u|� �>u$�e$��U6���><��I	J���ڂ��?��>b�	�H����\�ne���(�4n�%ȸ�7�dWIqXc��>x�ق��	&���m�K3m��K��{��>R&@�mQ�f��_L�j8t�X u��o���2�M�bip��*g	�lJ��Sp�W֣AE�M�xBrG�qz���~a;��'��LEi�
�-D.����%���	�P/�p��SYfVVMօ�Фp�&�(X��Fb���{?��qA_���̄��ÜVM���뵉}{]<�sƓ�V&*�1�tӺ>�\����d��
��`���lN�5^b����;(� }�U�*ń��yFcR�!��:ʤ��4������u�9������/=H7�`�g:�l����o�w��7�!�C� �e�[w�Jͽ����g4A�0Z]ӧC�CDș�@韂s};�j晒��
��9�
�ڢpC�����t҂�侯0 TK�tg��RJRt�ؖ�K����"wpZ���)g��X��@��Ő!�0H�g�Q0
�r?m����ʸ��3�e�/��~�~0o ��3!H�@� �� N��Cl-V�j�h��`����2D�Ӻ�6��~b���DӞ��f=Q��>�ā��`"W�Q1��GP����Q^A0ژ2$֏d���G���N��Kr~.R�v�QuR 61y@��l?��V϶���?t�ћLc�k��J6�Rj&[0t]o����LgW� h�q�<����A���&�X"��zE��q�S�Q�޹FH��&��;��=�\��+����Rz��Ȱ@��
��[��)k��r�~�Dg7�x�9Vt�z����51�'9�꼐�Cu��7c�]_7�}�dN��W�]��?d��b=�ũQ�&l 6��";��}�����V4�sw�qָFױ]"�4|�*a��A�l�[pH�]�n��K0v�&j�ޟ�d^W{�<���FEm��ٮ�k���;��&��������	�}���HAc@4��W�`��led�PR�4�Or��b�%V,�	6���)T՗���*n�لߵ�ּ.nĭ��<7`��of�+gtK�œ_��坥�	N�Dq2j6�Z$�r��"d�[q�<ߣt�2� M�?Chd(X�D�;��"�?2�a|��W��$��SZ�orӠ��4��(�U6�(�n,�P5=�G� �d������t">Cd>����E�^䞨�}��*�o�@5����Lʥ̆�l��M%���ސ���*���OsJl�u���`pE�D��/��?�||z����+�f����PPYx��E6�'��wq)a�l�fy���W7�.�<����B	�)���x�lUѹ��ͽd��o�H���DW/��;t���(�k�J)��ؙ؛�GP�G�2��s�h�r<r�g�cm��������oGP&g�-�ٷ��S��|<ϗ>�͕J�A����it�G��2�Lۗ��F�a&x�wk}/��y�	��GQ��g�?x^a�x��F��C�l��-W���~"ڋ����6���k�����m�@e�B�����f;�O
�G�:Af3��t�,�?�[�Y�6]������b�����ֺc�<�7t��0>Q_�.�|�]ae�,q��������t�_��,_��PRla#q7N�a�ѫyk�[���@ɲr�����HEu�)&��pƋ��hn�ΊrC�uB�/��C�.���a��Ɯ
�cAxQ�"����8�y�-�*ʫ��r9
^d&�5%:q��k0x���^\kgu�[��d ^ԖH�nO�Z���F��7�>`�uJ4r�~[�:�fsՋ�$�{�oX�#@����;��e+�x)�����]se;[��E�+�5���Qz���H������;S��a�LvT��57��nOd<��ܼQ�b��%�� ��
"D�����k�R���Y�����F�� ]�'�YD�D��,�m6Ox����Hp?�Q����{k��֗"�t��G@s �B���I�	 ��5�#&������K����Yt��5u� V~A)���.gK�j�}S&s�׽l�eO4�mt�("	|v��^��^>F{M��� ��#|"즨Η{��#O<�����M��~���_TrB�$yʱ>��5��O��i�5������r�c��Z�<պ�[W�v?gVͅ��f�3^Hb�V�!u���I�
�T��L8�T��y���/r*(؊�6PU!�x����<��j0�|>�;,D;d�[l�������H���WK��\|�������@��ȍ��F�jn ?$z׏/%
����-7I�L��U+|�Q���o��rޜQ��O��8��.��S�P��B�/ҷr͐"�dN�8�N��|:�ȣ�zx��;g������8�#I_����\|��og�(8f�N���ˬ��o�0��D�k�O6&��쟛�tn���z���sH������ u��A�!vԀ��5�B��&�D��h���O�Md��,�=g��讅�65k̖>�C��蚹��,�T�:����-(/(���/�ƾ�E����#&��2�����s���4��'�\<��2b��<�S� �<V*��n�HOs��c������q�N�
1�B������dƕm.g�˱<T��Y���	�����O���ȉ�v��SaW�*.�ԗOי�xP�EcO�{�s����Ub�~�pG��p.����������.Ts�1�Lj��qyJ��.�<��杌�+R��]���q�J����l�쵧M�j&���������	c Ԟ4I�s�������
����+���q�j^.��K�����6|�(��4*�ƘQE}�e�|-��0�j��:۬�e����1]�ʻn���}I��s[��М�]d�k���!�x�ϑ눲�W�\X�[WT�N[b����>oct0�(�)%�m�.1j��'��P�Y�j�;_�A��u1�0�z(�.&N�>���`ޘ*��L=u���]m5��4^�r �xf�v7�}�XVY@0�3<%������t�٫�_��a��7V���":�_�r�azn�T���U[�yS�ǡ��C��_�Dr\~J�58M>~�����WI!&��/Ov�^���a��U��S�_H��!/���{�=�V�����	��0��<�����R;�\���O�|��-fLo�ܨ� �:�䫸��P)���|7��)ð������>8��b�v�~`��z`J���B&-U����t�`�����ˋ
���ƈ��ù{@5�m��Q�.�� B�H=�J���5��{	�tA�t��Q�^�K���sO������H���Z;�{�Y�9�\x��`)8QTɰo��ދ��*�_PY��&4!+�-���KNaSy �[0Q�`=�!9���D�TY�������سn/n@+���������
�b�w.��4p�j�W�]吅$� ����Y��܄��RZ<%P�H�7�
���
�"�GV;.��f��k�Q)�\������"���^�s&8�!�@�,���k@����w _�en���R���B��{�yj���2�n>�����<��]�zHٯ�c�Z� M9AHCX70=p�LBCK?ŝ�xV:���^�PC[5�,�k���P�y@?L*����,0!�m��rk�
�T��BGX�|<�	��O/�j�3�qQ@���ߐ�#�8�L���_�/~��{O���e>jA\5^?EBi������,�ׯ��Ñi��]&�5|ߑ�v��q"mBI0t�9@��(��n0�5��_b+��('��O��@�P4�5S\k��(%it����8���=�c�1��B�N_����d�u3dдWe�@8�oB��34�(4�ӿ1�bo=�����[1�EÒS��q{�5��Q��<�E�6��@������T|��d�M4!�#!�1j��m��m��H��#�n�2ms�P�u�D�ϋ*cRslL������[�8P:��K�~W����B]k��efʜn����_�&�Tw][y�.��>�پ]��m���>�_�2�����Zvb^�.f�U�hD�4^磚��r�>���M�H>�g�n���r�xOO��˭�-c��J.ZB����cS�I!]8H�{��M{�g��h�����06t��dvK��BJ��ػ6��r4�/�����};ǁ�u��'�-˒����e�|��Uu(A��Џ�g]��ag��؃���ٚ,�}�����¡��]�[�A-<�0J�����7�
6+p�&=?L��7�H�ӻ��Q�3�A�dx*��s�lD�z#�	9R>�I��]��\����>O��Jvu5�P`��x�k��UgERA&Г����8�V�"�C]>��(��{��tY0K�qx�9�Njs�ڤơk^��y(<�:�
�s�anK��ˎ�j+����M;U���f��y/o:]�xaq����pg�i�jU�l_Ќ3L��L8T���.���A�!�{����I����H1�;�25+o�*RC�K�Pτ�C* Q��T[.�n��?��^�"�'�e�������3�ķn��T[�D{�+Kcc·4,�L1�R
砪Z%«�Ó\�z�>z�{Y�Ԏp~w���o5}#G.��ii݉��"rQ�w0�j����8Xe�y��6�	DD ����7N��+�+O}��5w\@+�%?�2hx-�\�D�e��m��p�h�Z^.�i/E��
7*���^6�~ܚ�W��#"�.6/��_|��&r������#߷
�dlk��r6��rd�1M���J��úg�]�����faW��ձ_5�f��Wi)��y��A(�pY�}�!1Nlv�3��Oh�J�J��eMeM��]���7u�7ci?��Vf�[�"\l�ӑ,h$	��fu�v�(�P�F�-�ͧA�d(��X�2� �+�l�L(Wթ���N�U^��O�o�t*u��@�(Q�b��P�0mR�mHw쬬���*0,Wǆ�>U._�wsE�W>��G:�j�P6�C"�{2Usq[m$����^�ψ- �c���u`-���0"������D�ldO���r9E��l>ii��y��ZKه՚*S�B�~���B"d��O���t��{%igm�?zW�oF48Њ_s+<�?�t�9�V���*��+��b�8-k��r��  ��8��"/WI'����RN"9��]�5p�-&f��g�^�'�Z��_%M�AL!>����7n
0�)� F��R�@������:f�y�Ea��c6�Ĩ{�m�~��c�Gw���$Mc�� v�4�u�����zWA� �-�!�Eޗ��OY����e��{:�?��-�^Rԃ�K9�q��|Em%朄s
�oƋʜ�Lfج@4�ᅁڼ���.������y��k+�4��I�?�Q���k�*��*���6�����H��5��a��`2�����Q��T�-:�ֲ�Sang(9n����A����H�T���v���o�:�7�:&ݰ":�1�U����n���������BG��;�{ả,z��Q���Q��N��uM��ߨ�����!��I�����j���z�?��k.IC�1q=����$�pTV�W��t2@�J�]�_�i���:��ʅ��\�`����xB�])G�nM�g� �r|�{�<� 4�?E��S-�p� ������դtiM}[F����w,.��n.��{�;�ǚ��(��o���
�	�
PǺ3�_�X�'���ԀckL߾J��5����u��P��~�)[ܣ!�ÐI�%�"��!͂X|�P�5�-犵�#�R_dŘ�Ŗ)�;�t�-`���qv�I���@b��Y���A�c:�`P>�`$K�\�.B�U�R�Ȳ�����uw��ATI�Ps�7ߣtr���|D2�(Q�c��?J��{�yHH�<���Ho[9�*ٯ�.��S�Qai'���Խ��X�8Dc-˒�l��mzNd7c���ϧF�[�����H�=����g�R�3q����DZᝯ�U�E�l��}�;BI��w���/��{�c�����M!R�@腀��5���I�����Ы���Hމ�ˏ>9C��bZ�wty	��wФʾ��R�~�r�N���b�7�=����R�E�^����.�=h�����΃�������-����{~��s�Ζo�5�:�'�P��������t�=�f��ۥH	�[J��*��[fZ}�5sn�{Dk�,D�p�:�=�Be�H��f�����{��O���6�n��w0�ȭxyi��>Я>�}��')���F2�;��Qt��KQZv<�Չy�p��?�������}�1�GiT�:���,�WK�����M����l�ۊ�WV�g5i9�N5��h�3pX�-A��K�%�9�H��C�O`o��w��Z�½���0-� ��Y�99w-�^�޻f ��ip�q7��n�1���9H�<�dwQaG6tk�VyM�Ű��i��yqt�Q5i�?bp_O�����elʈ��K�m�\���s�R�|`w��|��gC���y���j���-G�s�'��m$�V�o�㍎;�\�Ճ��3�RJ�ؤ�,/�GU7:$^�������-c>I�h�6P�(i�˺��8��N0�>�B�۔�6�!�}f��R������LQ�[��� �uK1ih�[![�֦��Pl�/^^��]�}�(���8�$:XԾ?̮.�/H^Wu��?�lF���F��ch�gl���O����P��uLl�⹊E?e~e��#`�]����.�T-���g0a�~;�UJ)�Q�q�O������*S�ć� U��ONQx�R���C��7�KU/�zt�U:d�q���ons�N��$ą�=-��U82�s�!��HN^�-�|�#��/�yT��C���,H�����|���b8ڷ�WS�,��*I��el�M�?c�����՟����{��Htָ]s�0_�ۊc8���UV�������x,�ǟ1ɏ��6�e����p�f�8i%i���_V���� ���麺�����*�P���>�ۖ,����F�U|��nTT�ϻV��,�<t��)j�B��������.(4�aMaiQ��{��)�Rs/����e���l��c~�{Nt���8�G�l泜\�]��p�J�p"GN!�9���uH�x�M*�r,zx�A���%E��*J~+��Z⚂����nّ&�1$�#
�H��B�2�Қ�o+ҭco�S�	m�k��%RƔ0��9����/�:�f�-�O4_�0�6;ʟ�~�L�*R�HE�r���r6~=����X������
����b^)���{��:�2�`n�-��԰���C�ʑd�_�D�=�՟��G��ݔa���'p�5萠y�jA��iy��Ė�C��~�&�{n���}Z��b�������b>�}�<\��KٛkE���&����ͧf&�����N�Th�d|-P`��3$��yic���y-�R�I�o.c�?)��a\b��:�����c�/�����P�ڷ�f+��i�*Wn
N f�,y"�6H\�.d9���ǉI.�.d��>�i��I�>�LE]�3���P���>	�s�������w�#�wqM��Щi�~)�I�]��F���}(m��aܴ��y+�H0��Ǆ���o�ݮt2�]�>˭F��O_�?�a��J{TNrG{��Qy�׀x��=���*�Ec����Ql�����|�A��J����kPa�����������L�N��ʢ8����9�A;��7�L/��2�UG�(��'�lP��f��A��F�Sgo��]�7;kA�J��J��d(�Z��f)q.��flgG"���޾GS_�ō>ue%�<xp-J����z�#쳎�_�}6C��VT�x@��^� �l����>ӫ�/��Y/J�-�˒�or�§�*��-�d�|��������h�B�&j��
S�RTH�1#V���Պ"��nƏ�vΖR��D:�'^�K ����ڵ�d>�!'��
�Mc߅��2��ȇO���:˶j��f�5QV��.��5.�݉�^����Q"L�RQ�U�<���qin�j�݇bF	ĭ9K(u�R�Šx����u�N�5 �"7�T�d.��ͮk�l�D����Ȇ����Z�i�;M���;��\���2�x}������Gt��Weh-�]��J��g�k����}�"�:�����$�-��W5^�M?���,���~]x��7t��v� ��|"�E1_��R�����fB/u�RdQ4O�h���^w���w�
��"�O� |��I���h�qL ���'�.���bJ�	��)3���L}��32��TUf3}��9N�O,$�)���(��X�s�o������\��h{�@���1�x���{C�J)4�b7��<[�$d�����C�*��Ƙl�����BHnW���v��Q=t�&�c|�}M���R��Q٣Ob(n��Pq�Gq�.� �`�N"ӘƋo�"n��s֢_����b�dy��6y��ԤR-=G]��2Q��4)���B�r���V�EC33�ʙXg'���iP�yIMrޖ-^����8���7��Q�zm����2�M���G���[w�R���J/U�VV���
�e9�7���/6}�Բ��m�f���7�6�<��-�k�fAB��B��)**�f],F�D^:��2�	�õE,����%���ܿ�m��2���c�FtUfրw�c (�]Y����[3.�%���h�qG@�ɱU�ܦǟLP�ב��Z}��W��dݏQ�`Oh$��3_qjB|:�Tp�^I���F�N��+�f��XvP�읈ƈ	FG_"*{���0�><�L�-�� EF�Q�<12 ��q�?�2��"OW]A�S5�]��z����X�
tG"=g���޾S`_��9$��)��qҧ�F��Y>����u��S�Kۂ�PY�|:��5 K�ݚ�~�
+f`w�+ئź#�5|��>4:��<�՚���V|)�i�݀�1Jj>%ٜ;5E�5� �~.M�O>�����$�d�Dͪ���V��(M��콣�/�c�1v~wx�O���{ݠ'�fv��lQ��%%J�E��֍�A7W;�x%�33�%�@�k{�3�^�L�tp��fu�5'B^�ӨנmE�B�-)%�%����9���ϔ���1v�#��=�!�Z�G����淀�S���鵧�
 x�^�� ���h���#<UG*]�,�T�3cu�r��������~t��%M�xoU�8�M�����r�����������0�mD��������W2�Te;�~Ү�A�{lzW�����߳=��a�R)�q��;�5��(O$X�
6�Dl��P��dFd�o�PJ��X
��M͆-�<NH�5m#��S��B|�%�ܢ#��b��Ԍ��K�`�h�Vl'w-
���Cay.��|�B�L��9�Z�˅�v����w4L>͋���l�	ac��R�6�3�U�Hwq]D���0�6�"��0��9pw*}x��V'�8�_%<���Ż��t���W���3��q�]X-�t�#�.U�F;�ܺ��U5��������ٶ�����u����ܵ�I��|M���晸t���G�i�q$�MP|ϴ�MT�#�Y��}#��`��%�q��>�Z�w`��(*ʲI~�������ȼ�e��Z�-���a�|������Č�����d���Sa��\�7oʒٛ&"n��{;X�A�+ύ?�_Z�Z�8|;�/���\������UEǽP+k�W(�Ӊ��̓�m�6;B�ҦC�@�iw
��,S_��9"sa��Tn���~�p�O���S'���>�(_�/d$��ɣo�:xw똴�H��&��_�b.�����Ik[2�N?2�{~<���f���|��i`��+�	o��OK�6���ָq8�2V����V���#O�:��V�+�����r�;.pK��K,�*�c3D5[���2T3)��b���|��˞�B�?��X��?`�;u�]��'9�Y6Ř!4Z	��`�S��M�ψ��k��+����SwA��*��X���C��W+�����uT^6����ט�l^;s��H���̪�d(��Q-�|�G��b"J��Ec[[:J�b��ʉ��o?u�R�a�̱j����� ��|�����k��K����"�4�N�c���'Z�Q�K���͞ͅn&�� ]a�����7���N�MDŮ��_�9�9�Cl���Xi�	��7�61�h�z2�Q������tA9E�we�?t�`rm��y9��(���Y�H�h�O	��vu�.��;�%������f�Y`a�������?�'�M�HM�D�/���i6�T���#�J��7W<�M!�(�6�1�5�c��K|i������g��&�u?�gV�=��Y��Z!`2�O��V����M�e�c�#���>��>3�$��k���*�9<$�N�B4� �k��v`��5 ���yhm���pn��� '����}���D`&e�s������m�SgQP��"8gT���nL��uE�rbom��s��}�a?�pS���W?յ�;��^���	�"$�È�!���7ʕ�s�֏jG���CL�v���]�_~�"i���U����iM�,�mb�j��TE����m�U1����m[��'4�$�Q�c+�ۋ��t��鬜�[H�PſPK���%_K��+uĢ0X�����=1e��qX�ȖD`"�DI����59�t)_W��kV�h�8�}�c��~S�̈́��e�J��������櫩=9&�qh��T6ud�!/�����@��WX��;t1�(��ji����p�:�N&G���@�;6�S Je+���Y���o;�Ȃ
 �1�_�[������*@���b���ޙ_�i>�bC��_l�r�M%N����[���لi۪f������O�����������A`�ׇ���Q�V5\9��_�5��ǡ{W��e�I>ǇAy>����Sm�;�s١���J�b����X�;�����48y7��|�����<�!O��k W�GTFm��jy�}�B_�Y�.�3�#ٛ
~\�
Z'���;�+]6�+]�H���c�=��h��To��.B�"	���p����B���G��[�����j3�>��3��j��=~-F&���,H�P�~)�N�X�>1��"�������Э��C��v3stt�T���o�'��hӏ����9����� �Yd�J�P�c
j7D#�I�K�>��'ԱB��|��kx��ƕKnN�)Ԟ�>٠�\nR`��	X �l&�Wl��r�����E9\m�z$��H
�5���g�z'���( �����X#_Z���#����k�l��>J�1@�w��&$��O���D����5�R&�'�2O7Q�$dN�F	_	p#�֘.%�����h��,u3
CW�������h?��'W�i�u`
�4�VR�s������ !�����Z;Өemq�;��\������&ʜ�v�L�P����gX���<�r��E�`�n�^�E���y�0d)zTe��`�7�s�\�_��o���-7�km�J��@^0��wnE?t���[p�:Z���1�eq��J��^H�V5�x�*xV���sg���sd��5Wǅo9�,���uҧ��n~�Y�ơLj����(eo�f>�>�s����C��b�q��/rA��,����%�WAz}�����Z�ZI����m'��d JoH��,�9�r������Ir���H��J5ePEC�/O磻{�U�Fo��5����d��=����eދ"{n��0r��4s�]P7�r�N��|b��N��ж���ցj����_C=��ƃ*P=����{ma30�~�|�g�'�P���~K$����Ji���L׼A�Eu�S���7�O�ר3�vp���|Q��3t(�ji)DW��6K���&�n,Գ}�w�<S<ww����Y>��t�亙 ����(\�Q:#J���05��f��{>�'������&r��)>�&`Na�ﳼ jȣ�o�Æb'�?<L�7DM����X����|�ԓ��F�f,%����5�[V�����@��L�g^.���\��b��,&��ȓ�
���8U[����ޕUmp�`mW`dV�n���F��DZ����<M��r��_Љ�5|b�`����+�����_��m�ȧTV,v�bb����>9�>i� ��N�%�%�rTf��V�7K�7�C�<#�{"c�t,{�>h��T��t�����ȥ!�s��|�}�p�m��1\�c}?"��d��`��gB�釃Ǧ����FS����.���[�g=-S�EGQ.���WU�#��`>��%YM��%:(��N�5�H�H>`�]^��LMo��~�݇�nD���+e�o}�K*:�΄�n�N촏��#,�{"0�l��X���ٻ�z���R
��)��=�߼\ b&������$7C":��4�|R��A��J�b�ap�*׫Sp�IX*�5m9-�f[�dD+A>D����x�1�[�	]Z\@�[�X���	$�,e�,�©��G�JĀ�PY�!�wfZ�ڽ%Ozx
��"���B�{�B��<���p�V��~�t�Z�E�>�2��G���]a{I*M�W̊�j�:&{��TX�u�d�G�߸Ռ��YZ-�$�ꬍE�Ui�����i�i��iF���٩���jn�*=Q�*�k�����Ԛ��w�U3 	�Q��� �Q�)��!J�m��:`�'�7���괁���ږT�}ne�0��I`�������=�8��?����8�����av$;�.A&j��ٳ4x|�Үڐǟ��ո��p�l���Ğe���'ͼ��ռ��v�n_{�����-u�B���"I����Z��ȣ�{�+��+��ӑs�w#�;9�f&8Ր��c?�x���ܕe�n*���>���P ]��V\�s����#	]���-A�b��ق�Y���o���� ��A(~$�X�E>��"��V��Y�Ԃ��bo��x�6o�2���:Q�.��Y�Y1}���oI��Z��!p�)���g����R������w�v,�ͺ"F��AEb�K���@6^7�N�d���@��Ҝ{cQ=�'�i3�^�嚱t�K��������V��o�C2n�F���DX����Ej����N6
��~��l�����7�>^��WK[VW���k���x{��ت�G*�5`�6��l�{�C�����~�ި���I�V	����н%��k@R:�|C�7��BC��0�潩�t;�_s�+�ɞ��*���<�pmʷ�*�8�Y��|s���~�V�ɪ�{|H,��G0�T��,H�/ו�N�Ǟ�)U��!��*X�I��6u����{�/�sʛs_�H?�]��C"��g7�yҠ���	�v�����ɉ^gms��(�Y'[��`tK{�p��ǋ��������L@ �뎺���B󀟛�FD��>��\�+�3:��S�p�A����l�߂~���5��)���,�i&0����M��٫ު��[��,r�]���Ҕd�39����S6��_��M]tc$Kķm�V�f'���Oa�N��uZID��Ѕ$v�cR%�$S�dơ4;/S������{��M����|Sg��Z�Pc���yߴ̘q&N�%����7��#J�5`�����-!�)��+ݕlO>������vO�iJ &�m���x��Y�A][MGt��~�C9�f�'-��ӦJ�N̶��dJ�8�T�T��y-fIax` �1�����=���G���Z?�_�w�=�� ��y6`l�1v_ax�Hk����̘:�z��5$x��hUn�n�sv���Zam1<9����ˎ����{�]�����_�ƵO�x�%~U2,��à���ꠉZ�S�o�V[�����R��_�jAo��{�3!d�ZL�h�(C`%����ۙ=�� �f��C7HT6x��ֺ�XejTT�U�S��h��,���V�˴�M��DGǔ�����2�1�v��O�4>;��K�*�w'Һ�l4�;q�AE�Z"0�8h�j���: ��� �x�R%����&��S��5@�E#�*?�sJ�C[9�='�͇�~|����<�if�4ɩ�/��7�S��(���fS:U�s���
�Ӗ>ܝ�C���HS<�g�sDq�@G_�L�!㤆���m�~�=ԡ��	��̍r5~�V鈳��Q��G�l�V���g�Sj`�s]��-��`]�1�%�}�My�;��Z��g+�w����O���S3� ��G=&����|M|�����{)�g,�j���|+�)��0cf����%��	чaWYW�����,_��&E�W� �����$�]��HXSp6I�܌�t�,�Z^����17Q�d83R�d7���
���,�'�X�,�w�V&5$�L|6Ve�]v�$�
tW��� �ߒ:(���2S�D/�Y�.2��b�Uօ~"�5�s3�p'�l�M L�Z�pV����Էy�<��R1abG9�(��t>A��Ɠ&V�/%8�+������ĔѪ����4&�j�&

������mS;���͏��e�թ�����4"�ec�K"s�_�y����1R���jo�[��;� �s�w�k|׻<��E���U���J�� ��QQ=V̋2I*�^M3��M�+0<�a��#c�g椴ʺ�����DM���-Oxd��\�_O��s�k�tv���X�s5d@$ؿcuR@^D�V��?T�Ybs�L�;�'+�H����4���J�scQ�Y�16��n�i"�R��p����;c,k��{Е��v�]E9e�me^2�k���궇�ެܲ�˼��'ix{օ�X�����D� "��bV7��5�_�9[7��'O@!o��S�ɹ���!"ߧ�k>�D�,���Q�qJ>U�\yN���՟��|K��0����h�%��)� %�)�'�L�}>t��V��".\wa�3�ӳ[�Y�{�Ks�}�"�y�%ǥ�=ʐwȫBb�Χ���qo�U¥сUS�٘�v=��M�/eBߊ���D��Dit��*�1$�R8�@j���J!��cʒ���8�m[���r�|�w:Մ���d�Z?
��\��I��D��'�� KI���vO� �#�
����!d�,��o&:����&$ru��M�q�pOF�eF1������DW�.�_&�'x���?�v��0b}�����f���M)�7jSk�M5�V�z��@U��Q��k���G�e��5��
lA���+/�����.(C"�Gqz5�4��.Gl+����_��� 7�d��Ǧ3;��w~��W�n�9��K��{��˾�V�I��?\�`��t�cG1IT��io!��v:$z\���p��&x�[H�fd�э|?�q+g#h� �c;�)��|����o��fj_f���[�nQ������&>S�_/�۳ܻ"8g��b#7�}��W�`�I1�>(�Y��M)��x��)�rH����z��6�o;��r�����:��E����]N� w���qڌ�A��wwTt]�-���D$!5����y�<��$�ѪP�O�E��j�n�i]�cE,�0��Z�=�<���=)�,V���l�At�QR������͚�K{�݅���9�w,~g������{%*'aG�jt�q;��R�����lt�K�_�]5!�aŃ���Y^6�>H��ք��M��ǩ���6��0�^�h͔���'S�ށ����|��x-0�۠��v��ձ9�āX4f_������x�.:G���T�R;&�;b��Q�ko������=$�}�$��������nlX��^�� ��9�Ľ��<����P?�n�[t�i$�Qx��S"�"	_�|©�̗sZ�\��f�;���$�+�s_r�?����g��+�� � �(H:�)��6e�`^���"��]�<��'#q8�A�z0��7�PEp��~m��� v�e��FOy�0Z�?�-V����&�؂�\���
�A���_ ��"��?C���w��MfYk0.I�qH��\1/z�z=��-��[�9ܺq���n�,4���C'��p[�O�9��W���;x����qT�f���d������F��Zg���]��0��A@s�Za�߸P�.�-��[��9�9^]W��A�-�2�27�(�a�*��OKM��2��M�IA&�Ba��.�JJ @�h~7l�U<�:9.�DL@(�q��Z��,�ynL������� ;k�w�[LDkqWB��g�p:�=RZtT��	,%+V�l��r	�����s����S�l]����I*�d�?�q �$9�C
��>ܨ��ll1],bY+���Kl$��[Q�`�f���<-�#>ۘ���VN�<:Oz����:�q�G���p����oj_�����>:<��d6T�8�҅W�xa�69��@�o��)*�D�����vW�\I��
%�D��PWB8a��b���ƒ�~���]hX`�&�N�c�'c�!JR5K�� ���x$������\�i<�T�+@��OF�"�i�
P�9���%���T��l�-��3r����V覺0�X�@���'L;����%��ӕ $�H�.��y2����ǋ+�[I�kz�3ղ�a���O��Y)���Q
(�A��PcU,�g�o�;��}�;/����1hC������{�R��� ����Z{Na>�V�c��W�߈:�Mܪ˵���`&1}�u���m�x�`*U�
{�آ�B�,ٞ����9^��-�@j��^��-=�_l���M��RR�����5�n��l��j(�=#�"j������ߦL��5���(v�����5Go/2>����h�9�Ӷl�r<���b�#/?�ҁ���W裏z1�H��9�ٳ�W��N�F��܂�����#N��M�43����e| ��^�o����[�#:�6��OG������_���^*�*&@�c�cX��W��訳�ù�S����.03���Y�[YD�酊^1t�iȶ�b��g���y���3�˚o����֛V�e��Nj��tt�9F?Hx�������\�0��O�s..'ɋ���Y���.��?	�Kz�t�X������L}�M&�����\ML���2�5��3�k ��`�w��R�/&��i����v����w���b�V�E#{l��a ���t����ɥc�]K����p�5����ʈƽ!��h�W�W+�Gi̽�S��
>�Aq���l	93�׈�Xg�4�he�G�4_	�:3�v��+��8e-��}���"���R#��Ŏ�,����@2K0Y���v0��Y}m�<LNm��p��4��#F�URR�JYi�lp�o*��n�~'���W���2g%Ř[��h�|H���Qi���ʌ����#� �W�X�+����[w�źT.	��jAZ��	5fT�-v�Y�>�
�UӸ�]o�4e�˗;ˇ/������|l��^�',쌼rFj@Y�=BX�_t��83a)��������,�QÛ?�eY[lQ�3��_��?�O�c�i�����wzgcF�fp���l�N�3F
��9���&N
;0n�A�G�/m����k�� ��}���k�t���
�څ��T[Ⱦ�@H�k�Qj�4/9��T��\0m���
��6ǐg-a`�A�Ui���e��ֈk���oj[Ӎ�E��Ecj����w�g]�Q�� "�P�����Vv�=׻|���n��fXr���-d�
�M���fχ��^]N��|�$�� A��5Ĩ��R����_|KG:�<�(O׿�1��!������	;e�*j����S0#aE&|5�{Q�]�����&�̴%���ip��xU*)��9�V�-�+t����ov�R}��~������)8�В��ʱ� %'[Fj�oV�i�b�M ��PA	�5�m��
n�Ŕ���Oط���˸��hH�ldH�A}z�e�G�˔fG_§��D���O�9-�H��0�ؠD�Ḡ�f��](M(���s�[2I2�k�v��` ��ە���4�۟���#���i��ʳ��%����.Jw5I5�a��5��\s�gA�������,e�;m�+t���4eA�>뎏�_{�ᶂ��2}�����|��	s�hr{��V��ݗ@`|Zs"�Y�a�-�a�AEXf�`H������g��� =���Ȗ<��~n�3�wH���f(��i�ŲR�a��5��}`Fv�_m�� ��j��n������i�KN�����I�8�bQ��\�:�-b�+3J�uId5�+��{/����&[�`�52���BRW5\����.x�*$�7�����m�sq�8=׷�Ӄ<�aKy����(eb��Q����mK�|�(�.O��	+�^m&U �>�}���ѿk��ە��ɋsə%���}`=���� 	���3�~9�Qm]��nH�\)��J4����|�N�?ޤ�����xTy���w��5op�u� �]�"�a�S�9]!]���h������R���'����Jw�b��]V'�W3O�y=�ϑp��~���$23����
qP`�N�C���Ts�|�{a��a�ž�������	o���P�*�����1�-{���uY��9���������?&�{���*�C�|=ܓ��X�X��h�M�u��
=zw�^�&}���b������[�}�b+�v��crS�d|(Nf�.�b��2)�.�Zk����nd�I�o�}L౮|~|��xa�����>��'^a+�d���)���F��o�M�Gx�L���gA^�a�1��a]��W��'D�̜\��Udc�*��1ɛ�
Z{�V~U��d����|����Ͳ\��KTZ(fCt�z;H��x�_�i9�w�z;�}Hv���$�>�"x%� ����Ւ\���ʇ\s��Ec��ԛx:R	�F44W,�8�-�_=�)��T�M����)CHOU��}��.�,�0�;�T�s��(\�GcR��<�3x(f�-|�y17h�-�c�9���vJ�u#x#k��7I^�D;�^����������oap���(�9�(�m������qo��s�$-p������3�(k�bA�R�4��� ��5���߯f�����!�gL����A�ٸ�^ �n���͛��LS�1Wԓ��G�!�YU��_3��hho7���=�*�>\3I�(;
��|M�%iv�;��g�LVl�5`�g�`���K�j����W�O��2�Pni����Mƫ>�r� �#3o�櫜r'y���,��])�Ed����Y�ڥֹ:��h"}�"�U+Iq_��]����'?���+�0'!���~�nX��K1�_�Mz�f{�?vh����	�Y��;Tg�=��-ԛ~!�D�s�k�?��k���v��ݔ�_b�S�b����1�YCV~����fEg�߷�P�'ďA7}�އ��/����o����i�s��u��E"�H��ҭ���-tגX�\=��sk���('e:�D�n)�JYM��!(r��	|z�����;:����"��r�� �!f�H�9�Lv��
�HTP�j��IX�xĜ@^�b4�pÛ�b�|�sF�̬��;�ū�; ��{�b���_�u��Eݡy��28_z��T�*����i閔a�H O]��L��%�fұ�sZ���:�̋��Q*��+-�����0kw+:��A-�G��gr�:�ܺ�mV�Y*�F���{B۷�޳��&J��5K�̕E��˧)��.l�#/Fю��q�\^�K�;�������
����N�o��!����-�7��������g!��ҟ�h1��}v�b��b	>]ƿ�9x��:n764O��{"�������2,���{�(߯}t@�[�����i�N)�;����VT�;��nE�<�'�������9k���Z��<�}?̽�����|�Öo"�豂QW�p�����+��n��3F���JB�����4�s� #0����hf9;�טm�~\�u7yW��5i��%_��G�}quhUe����w�&�CŇ,�M��f'ī�"�*19��C1ã�t�ʔ�^��i�7a�V�1��w�U�C���)=����u��6���(Lj����h����)��U��EY1<����.%�(A܂(\1��걐ҳ��E�����\6��'f�Ӕ' ��A����^��(\��)<� �O*�N��tں:��{���{]��P���I�Q����sy��4�n�~AU����ra#���OU��e���J?���K{Ӫ��:	v(XZ�(b1��p��K`9�d�N{����S�ҩ�E����mB0�Z7hgۈ3��݌1��S�dVzp�X�n5���8������N�2V`m%!y��c$�hM�p��X3�D�]���8kϽ]g��A%��'ٯ�.07�5�v����N��]���H��G���P]^#��0�q���U9��Yg,��y����)%�߸�=eI�+���2T��K�9��g�@��[�I�L�@�Ss�.n�L
���_�����]Q��H����O�2u�oN%j���K�
�TU�Y���vc�?:n2��~���	�8e[,��j�;�c��xy�F	�ó���[ ��?lv�z��: ]bG�C���ؑu� D��@���m%f��	�����v��bN�`lCA�fV�k���GJ��L:/�P~9Kh/\%��h���GJ:I.�S�)S�` ��n\�A�;h��0ϫ�cݰ���rܻ��Y��i�_p�	$q�޿�;�(Y�N���B�����8���B���dͬ�[@�鳈"�wn���qE�'s��qn1ŧ*���CU����C��I�\�0b��fbj7U�:x8C�������X�`NB�x���G֗l�Ͳ�dȧ��x�p��2{�)�"<��ь�(�)������5�嵢N*���N\�G��хܫ�Jo�tD
����߬��9�3�׾/H9P����q����D�[�-`eI�����K��%øc�I�m���]u��G6�=J}x������${��.Y�l�|���km�/� ��)�-�_��������0�|�Tx���5VV3�5zI���"����H�i.{�5�=�3dEokb�I�&��c��XTV:y��y}bI�29Q�n��*��C�(�V��υC��UϒlXHѣ��ȧ=�����j]�C4��S�'sDy���B����W��|.#f��(������p�_��cۖ�]A�(Y(���l�}rb�uxXۦ��2rV�;t�_^�����_r�W�L���9�Ϧy�X����y����HA-Wܷ�/�hZ���۾���3���0>�ؔY�kበW��s�d㯬�����Tvdf���^��)�\��~�%;��G0�=qg(����*�l�s�T|pc)}&R�	JC'�����?g�n�	��Ƥ���_�|{oh����S�j���f���Y�e�w�=��wZ���-Y����|���:��������oT�~��=�������[�X�<�L�	�9r�_R=��)�6�Ѷ���B�|Gə{��*n"y�!�^J�IYb�|���Xf?T�К�/~��W�L���J��#|��9ନ�dE$nFDnh4�i�v��1�V^OP[���7Ά��z��*ks�gX���=�h5�P��Fݛ(��f��J:���s�"��t#49yI���c{H��I�q����+DybEwX4��ڳ'�[TI):��dV�e�[0{tm�j*��b�d�or���L�8ś)��w�L�v��T�1�Q4'P"��u?�Vp�k
���0�gg{4�w,<|��U�O� 	�T��~F QM��u�k��|�E�)��8̛h���(.�4��֘���&��]M��␃��X��8���dX zz	%�]�4OU�ʪ$[z0�A�P�:�{am�3�����"2���XS]s�1�sk���d{#-'��pc	����ð\v�����Dm^�˺V���v�g�<=Ib��	dE��ת�4�DE�������� AbA���� iST�ڱ�}/����J4�k�Dji�UTLU����d�*lFESOY��p�Mp8奠h?����z}�iC&�%"V*��J��L@�dE�V�i�R�tG7o�kBuv������e1��Vp���;
1�`&��m�2~�XeO<ǒ�f�Nߘ�R��O��;���ءf� �!Ef���,��T��w�F���W�fwC�4�X�&�؅R5Ľg5�Gs��N��s; ������3Q��\=�"z��cώʅ�ٸ�.�c\ ���HH���  8 �\>W<|j^m��RZn	��:fH��k	��5�u͉���-����?a��VO߱�=�;L��5�T����=vHr�"7E�,߄��:����#����"�{�h�<��=���
��U=� ���͌���\"|X�̫s�7d
mi�U��y/���*/�?�N�w�sy�3,2��/6�f�4������Z���j�S��� "c�����p�S�f���!�m�t�U�;���jf������-��;hC�\ѐb�I�aQ����q|E&3y"�Q�D
N�D��\^�T���Mf���<T�|���K8C"%�v�K.�)J��6~�+�7*6��̌��>\�
g0�	�b�7�d?���@�%)�{�C�?,�F�إ��\�+x���hi[(JF���0-$�������=�/u�n�&�/��6�3ا3[�}��� j��V���n���b�1���M�@��"�-9<h>g4�gf'���G#�Ⱥ�Γ���X�M1A���*~<<q]Ƅ�-� �*��eK�t��&d��A �+��6�Z$��[:ݏ�K�o<�G��P�Y��=�b��<Ud����/\��]���<�Ab	���[�T}i�$m�E�w5/��ƿ^�ˇ&%�՟b',�Vq�h_A�m�����S��C8�lo��)(�?� C�v�$��~'��Ů���ėr�8��}�Aiѧ�ćh�:�C�1&��Q�~����Zٷ�Vl�D�Q�H5�(��"p��ܜ���c�K��-*]�T�٥_ankB|d���Z�{T����*��{LR�����|��e0F��j�[&:9��s��󖢷 ��O[L�15�d����m�v��Ã�B��玪|o�`� �eYP:�'��&��T��$���6RQ c��}2���Jd#ϣ�I���(�kY��:�B�r���D����(���rY9�<TS�b��	��@�N�$��2W�_�jUS�Z����a�+�*kL�j<�H�y���,�H��?K7u���!��x}�g����5�>�SH��l7J�i��؅%i��`�rc���&����ȱtgfW�Ɖ�Q�y`}(ʰ�Pf��Q���
o��g/)KRŏV��GO���S��BlcW����3eה�F�U������R��#��ym�'(@3tY¹{�>�tW#x�)!	��8|��N�����@�NN
��q��I$��V���=�'zzznzO؟{�PR�V��>b�R.hW^^р��%�Ǔ7ŏ�հ$��|ê�.PG �3&��?�.�0�͆�G�+L9|��}�_�uB����)d���h�dENY��J m�PR����$��e.}����)=F��։<�ű:�HQY�߶]&@A�/S����u��Qu�VW]�\���� "�U���ô��`����%�����.�i�O���Y���	����J޾�JƜ��ѷ��^����"r����q�a�.��%V�!��S�˱SW���1�q=fٗ�X1�"[�ҹ��'a6c3k�/�rش�\�n�&�Y�$��2l�$e�_�� ��ߤ~}pz��.�L�y{d���M�u��\ щ!�׋��{{�p˷���^��l�GSFP��=;F��Vs���ˍEr��jy D�q���Z젍�����=wX>{d/��1������`��.2�+�m7���]{�ɯW���Bᦊ��fj&��Z�*���M�_l�)�'D�C{]��ίn���T�6���8��6$X��/�a�i-�|P���ݫ_�(��Q����h�1���/��W�xZ���wd��jL5���&�c��b[Ӏ건��12�ͻ �<*������)�[��M�6�+4�2�^\�t��M]yQV�*s���[u�#���u8�ʆ�d?O4H�Q�觿�������K�9 ��C!8|E�oZ��ބ�i:u>�Kg�B����-�)Q^ؐ���0DMI[*P�
Y��U<��E$C��e>��E�V�\+�ʷ�I�W3�.�M#�lr�
�;�j�D͢�͢:�R#��k~6�A����'`�8UQ�$��!{����:x.�UdA��P\���+N��'�d.
��&lu�)�Ş&�Iߺ��mdү������q�*�|p��b^w�`Y�E�D�p�i3���	Y�5�ʶor���,�+��k;�=6-���jd�#���*����o���e��e�� {�ڿ �
��ﱫd���i���+�gV�s'O�]���jg��z���^�-��9����4U��
�<RCTj9�޾{�$��5�㷇?��<���������ogT)�:�A^�t���p���6�d<���*�V���ml'W͵W�7Y_T�2��;�O��ţ�@y�QqNCgGeE��3D)��'La�=�Q�98�ԇM@kOC@�ƫRUH���*9]�)w�kmٞ��H�;Շ�V�� �E�%������Dv����>�� �o2_��J�X��6�ٮ_8��t��-�V=�\
"������P�(���Px��d�Է.��
��P�6�K����/��a������`8�u�r '�.��Z�#�e ^}�Q���d���ši��IԱ\I���[���%��%�P�y��K�ܭn�/m��C��ҷ�k��{�Y*s������D��,���E	���wBv=�H�A��݋>�(�/���*Lbo�Rڟ�J��|mQ�O����,��P����H@�y�h�5Y/1SY�8C��h�6�L2yZ�"�uȁ���H����/��X�rf:��@DW���QW�J�>�'��k����PE�Nİ��B�ee�}6�O��*|T�P��r��c�x<�q��>�
���_vW✜���Z����,9?��_���=k�� �ѽ.wL���r/OQqD��%��s�e�<U�c+4�6���c��������t�4�u�x�s]o����+R��>�c�`3�;�4GO1k�89><8v�.����ܘ��G�l�Q�>�n'f��q-�N��%�<�iN�+ܼNt�C�(MN�lp3�����#%�<�]���#bE���R��[���g�j��%�AAu[�Sr�/�5������C� w��1ۣ����g+%T������3/�v{��<��=\_g��݁:X;��ڛ�u��>v5�D䐤��0���X�vQ��(���#��X���wJ�s"_EAv]�o�w���oE���/��̽�d��e*�d+����y15��8��Z��/��
AX+�g=�$�_�������3�^��|
�Ls�xq��ҏ�L-tТ���:��GN��`G���7��Y���s�k��ϐ}(q|�e�đs���ʚ^(��4�	�n���)w�ҋ�i�ߧ�Y|J$��"|V~�a�����R�H�jP�+ p�(�):A�ֲ�y�y��ʕWv$�l��v䅈�b�ɲ�k=tV{���0�̞��F\�����:��{�!�59��/�B�����M}K8g�m'�vhۋ�h�7������A�&?�����
9��c�{���uB�K~�9�,܃M�]�r�M�`�އ�X4d�/���V���������(�z"(�=�1坝�΋o��!F��I���z�Q��e�2�4 $�L�$��[����F�P͐�d�ݲ�Z���� �6��@P���i�TnR�sD��uhtV0�)ǾoL��E���,s��`�/$XV���e-v81�+�t��G�rB�m'2LOr4��t�WU����X>���7TZ�u�Y+ܡW)��E�F��I0�%�˃���D�	��[@���~߁R=�|]�jX|�/��{J�{$��9ev�{.�I�N/�S8uw�5�b(?��c?��/�����2ٝ�"�'|O��!��1����'O��7�x_�eŻ<��|�Q�%���YUVe���w��ʳ-��>��hJ�s6���M;n��*el&�d�X�n�i�G@N���O�-�肦L�s/�
�'x�� /ٺ�763�F��[��r�	��c�#mG\lה�����I1�c�{���nRʜ�bu�XX}h�}����=�#.}���?u��a�֬0�VJ��+a�:��ړ6(Y����MX��:X�#ļzZs�i�η��)�恒pH��Tt��zY`�hU^m�[uG���c}�x�Jux�0R�oQsS'���bn�>���_?��⇦O��{�0��k��T ���'t`(r���a��!,j*��}��ۿ�3F�#���4<8!a��P)�w��8�L�C����2���>D!\͊ޛjq|I��&ʫ���5g�v�ȁ'*�@]�AF�s�f�z���?�DASv4����raP��,<�Edմ�p }>Z:jU�x-��AQ��7gm��b�W��A؊E���:e
��͌)�Ǥ��睈�g떽6��=dp�9��}����[��?����l����1����%U֗7�k�-��d	i���Ka+J��e�,�\*`���4@�a�Hx��?��X�o_�}������µ���c���c���J�)���۸���4/j�Ҳ���0,<*����j�gz�c~V�r�ņ����F�B��"�D����F�ҦVU��\u3�c�s*v��R��z%���*Y�8sC��ș�o,��-��U�Y��M��O�4�,]�Z��#�n����Y%�Y��}�,l>�{ɦ+��@X�YY�^B�F�n��Z���*�C����V���~g��2�o�C� ������`�x��N�l�[q��,b;\��G������N��.�K􌾐�[�(�6�}�����?H�aI�������և�!���(H3ӛ��(���b�_l�~����#8T:�ם�wQ�/�Kp�(�>t5��o�^3�Au!d�pQ7����>~�߽�62s9�x%G��6`�s�|�������*"�˓V��*C��� �N����w�$��ZJA�5SN��(�۫r�^f5!L���x$8���)FP�ҏ�h�Dɚ���f���u`h�`ɔ!g$�~n��]}/�SK���}��M�>����;�ck�92+��˱[Ox;�-/c��&|3��m�r&��tų(lOh	dvs4h]8*���Z$�m4FK;��H�_$�b��Jq� M	��F�Z�P��ITz����@�"r�{o�\��62����%���NE߹�$��¹y�v6���rG�hhQ'��ֿJ�+LE>��j}ɏ�P�4��䉼<S,#���?*97QA�/(2�ԯ��mܶR膙e�|��NE��S�)�B�3�{�.U�?��s�a27D���
i����2���Nf��]K�`%�{#������_�֟j��8Ĕ�7��˫���g܅aE���p��Y�?Qww#��V��m��x�b��-�e����-`����-�[�Q��U�";_8����:{
m���n��#NB�ڠ��!0�w`jaF�x��A�4����J흕��>�����a��ֱB�3��Ί$E��ci���`���a��/'w�.�Ϥƻ��瓙->�;"���/�b3d��<rR�И=������$q��/t�@�婇p��J��C�T�i���&z�ʁh0W�Ɗ�ᮥc���Kl��E�	q�ml2�?v�#��va����>�7��o����6��5Ӂ�7�`� 9�5%�!�����:��Eio���/�?,-0�7�s��Pd�U��m��lF��t{|�w����A�Y���<!�� ��"��m��^�Kcp+��*���W��}JY�e�G�B��~w2(��#+Ǆ�XSbz�$��DFX)����A(�,�����n8Ɛ�e~m1A��N�.q��*F���e�����=�X#��6�΀���6�fr� �Z�~�C/� �7GԕW%N�+	���\ؐ~�使sAcK����2l�Ǽ���u���tNA,M|*Q�J�opX����[��`�O�5%��Z��S�Fj��^��ݢ�(��)���Y�2�l���u³^V WO��
.C��H6�M��5ɚ���s���`s�ȼҜ�Ws�R��iX���4�O(j�Jb��7j� vS����\/9��N\��Wz�YQ*υ"nQz�F�0f��	tU�� %(�|��y ]�*�����o�|�G����#=�>0˾���6|*��Aƴ�/3=�B����B�T�M���IWh����_�|��|L{0 g�r�@|�Vq�w�<3���*v��kyyEʟ���M����lڦO�Xب�L���82z4ͩ��X��sF��~���U���ـ��{�b�1bh��)F(�YpZ�v�����-�X�U�[�!���L�R�!{��QD�������y-��"ؐI����P#s/[�y���{�==n��_�q	k��:��|Xre�PG�O�[BW��P�r�N�0Z�һ��[��^m�L
O��}�^�3E_2�H\�a�v���(x��!�dE���*w�S6ݸ�*mI���	�g�܊��
[�eT��� �s�ӻ�+<�H�����$���QPX�{8%�)^��$N�.��%�p=�Z�i᥉�3�M�]B�,|��ݗ6���)W�U4�eƖ��~E�9:�xo�d�'ʻ-����Ւ�A���z����3��-\�n:�_4<'�9�F�nI��7��Z��}�`��C����4���`�8~���#&����Ԏir�/�g���UO�����+-P��ށ���ޭ�ä{g޶e�޾)9����_����q?=��n҂0���u�Z,HC��R���y����x�iXK��zb}��j�qr������cn0��K=�9~��f%�>�!>S�5gWw�P�'�6���e����R�a�%��T��#�g~��"T��i��Y}Z��$j]8 7Kvk�Sr��.����I�Q���.�(��N����1$:XkH�M��֞1��O	ð�֚e+f<~��Q7b�,�[P��X͕��5�-�j%��!b�����9�gAI&����鎊�$'���Y�C�Vű��?Hκ)�_�ҋo����R�r=6�c�1�����ߟPv���\�[hb�����68]p���M���n�\����� j��o��R-	�p����۽[�R��>����$z�Ύ���Vha|P��7��Qr��dB߾Uy�Kɰz�M`���R9둜q�7��Bp���e�8�+������M}�qkA-�PS��H�M��\O�֒���s�ˍF���_T��|C��R���цi�'��; ����B���e��k;"�ģt!�s`H&䲌]��W>�˃�)�%���W�3�y�rƤ�(Ya$�g��D�1 W Z� "�N^LG:T{nЫ���/�s�[q|��r :=�z8aq�u���oN�qX+�/y�b�x�r*t~�y�'�O�7�eC~j(��?B�Ȑ���soc!��hE�('a���,+���n3�������TǄ*�%�k����Y�؈m�]�ScNu�'��_1��idNp�#Z�o�d8�6G�޷��{��;�kM*D�� ���?wɳӿa7^��g�Pm��I�m�t��U��1�1���c_"��9��jG�=�z��R�z���������7���_�I]X�|϶���V���AFo[��Em\iL?R=0�������"[����4l��x�:�����dX-�̪�V��,�l)�����:t\>ߐ}�O���L%2u�)@~����ʑ��h������ nC�0e��0�:M!�_w�uQ��9�C��1���������>�m�%Z!t�9�$ә�2��7���zw�D������7�7�ȼ���e�-ZE��c���W����v�)H�Zk�6�R��`9�Li�i�&�n�ظD�$$�9�q/؈�Q���_����ʣ�i��;M�HH$��z��J��=��t,0=4<w���:���}y���6׷�=��>�AB��y���l03'K1�mr�R=�����ѽ	'�g��d��ޗ���J�®_#:l9��5�J7.R�x:l���R�Q��)9�	�vZm�<��x�f2� [+l�7���G�8
q~�le�usV[�Z��s�kR?��mM��C#�����'��%Uf0��m���u��9B�ơC��aM��x��?�E�߰FD �ZE�ڧvNEUjS��ɇ�b�Ё1 �]��Ic�Y�����s��q� �E"w��gM��=�O�ۍa�`�vEٞ��(�ڛ�P��*8���gL	�� ��ɩ�k����iK��A:4�PG��Zߦ`�W�:��p�5���]��ӥ�J[�gv�d�D6�����Kndخ������o�-H�q��mh|�v?1.LR�x����ǧ��=|kn,��Q���-q˺������������˩���f�s�eI�9��iԔƌm4��� �r��u0�A�Qʀ*�_���WƔV�'9�Z��(0}64���f��D�u$���(f��h��m@ @�CFC@Dx ��� ��O��8��<|�x�4ܼ�Z�n���h4uܥ�����1G����̯�x�Wp 8IxD3�M�A�|%�]�|��§2��GPt+�	_x=��<0�kY]m<�<ߐ��;������H-�Z_7��jwH�g;n"\��㚖X�ٰ��ڢ�zh�,!��:���!V��]��ZG������)�L�4�s���
| 6�A�)*D�Yr�x�f۝�{�y;��ݱ�du�aV%˔�n�N�cQ_W�\���PU2_*��r�H��Ț7`횰f(6m�#ʗ�SGh%�a*1@�	կ\p�L�wE\V�gM�a��o'�u\צI_���Q}���v�x�4a��?}�n��b�Ȁʚ(�T^�J�	���wȥ���Z�t�	?�ˍ���I�C���e�EA��>b�ƻ���"��O�����ɒ�,8�}����xx!�[��� s�q�!c��%؟=~�uQ{l�o���ه��Ӕ$�g�El�Z��iU�_IK�����\���:+�1"��<=D��$�+��������暄��"d��� A~K�xӛg��E}Z��,Y)]M�*�f�7�E�[4^٘I}r�y"�8���3w%ڨ���J�q*��˳KY:�qn�!Q��A,�L�$]m*+.(���P�8��[~��gX����xL#�8	7e���g�L3Eco�h_��0��3[�u*މl����8�Q9Z��|Xe W��rڙ�F�����K8�`���z/�R�^3���(3�G0�|���Py��z���v��.�-��ɸ(������Nq�Zx���9�xw�S?�����*����l����;o�x�����	��i����^��s���������h�+�}���&`�W�hs,h�cQ�|:�k�_�B2���� o�A��""ǋ&Z~R*��Q�5O&�yM�P���|D�h_�ʍ��"�'����/U�������p\:���#����i�$�e����I�̪vyPЪF�X-Ӱ�I)���2\������\+p�%�YJ|A;��M �)e	��1>��v�w��l�3z�����[�Ŏ7�,�L�Dކ!#G
�u����]H�H-ג@l���+^f��R�ĴxYy�«T5T��~cRRs=��3'�\|�n;[�}�J�i�	!�p�����*H�<��ls�w%�I������R5��M��{y6h$�.�Y�6l$=.y�=U|�s��yw4���@k0�g�v̚@�yF��2�Y�+��p��	\���].9���Y��y�_�/�#�{��{*P��x����Qrh�w78^�����y�q��$isMP�\�0���Y�5�ǭ�	��ى2�S�U,��S���ɠ�;�X4�]*���-� +��tx�ꫫ�2@��K,�JൢJM���Yv�|?t�f(񽒇�M{��7�x=L�"�c 6��k����w��Ѫ?���X|�
ڑ��������5�GY�3��i��0\G��.�-�٘�����u%����
��*�;���Ǘ���k�B�2��q�t�(��f�6���KI&<�d����f��#e��ڿ%З�h�%��B�h���n0�8EQ˽I+u����f��O��g��,��O��6��{X:�'4Ff�������7�������0QЕ&z�t�	�}D����*�	���λ�Pr�4����@L4^��#�T�3I�w$�������9a]�m�l\/���H��Jj�6Ny����7�����R���w�}�U�z��\c|$A��f(5V4f!z�%HՁ;��O� ��l�i^ɆPF�Z���Ր�mm��*뉩��5��F�T��s-
-�ș�AY����'��r�� Q^ą��Xwy�g���8������_�q�0��zM<,+=�4P~5
7Kg�C>B�i�w� 7i�=���8�Z�j��X*���$��� �������/��]���֖��d�(琖Z{8��{Qٔ�YyS̓�z��-�_DMN)�#bYB�~G �R��s��"�O��P%�yi4���,3����d�.m���&����w=i�ӧ�W�p
��2N���⩵~Th�C�Z'�"G@�bt�����^:�һ�I�Z$,4��<%���@�NW\�n�E�e�"�:ւ<�e0��_r��ۚ��l��y�f]8�p�d��g"E(�-�{r��mꗅC<�]�r���}�J�"�o䢓I���M<�"�DK�~\ǡ�����O��򙻷���ų��h1&+�;Y)֕�i��t�.���=��J��S�i�s+��"�­OyL�mP�V���Ng{2)�T=:똏 9-&�9���PP�\Ȅ,�,��.�d���ev1}�Z��g���Nr�;�DJFsp�G��Z�?n�T<<�ycI���l<]�ll��fP�9*��e��e�}�p̀R�b��@��B{6N�8�J�<eY��O�E�����jA�^1͆9h�t$����@�e ͺ�4{�k��u��`VL����pY���~J��>ZG*��ƛ̬�����T�%V�J�K@Ų�D�מ�����}X������[Qdߤ�i������7p㔳��o�Q����"RZ!��K�*1-��1J���ʨg��㕦���GH� ����Z�I��S�0��Ae�?O���M��<��A�U�Pzc�$T�@ŕ��HYB�j�/�����u�%2~d�>֤�Z��R�)��}���v�F�V�S�t�7�O��M���V��N��9�����XMq�b�&���2��T���p>S�܎�蛇G7+U4�c6(D���&}QD��H��5ʹ���jI(7����i�+�T����fy(�_%��/��~�_Mbଅ�L��֭�>��u�)�ԥ����.�"��a���>�Ġ��$}�A]�I��a?O��A�cB�)q�+�$g�����о�z�(O9+1K�5����v��}�i�������'��;�y�⭒��I�0�--�y������Y�I�Jf��`T3��`��!aʒ�P]��Y��>R�K��X|������!����Bj�Gx?ʰ늍�sg��2���Zg>�z@��5�Fכ<&�c����(��TbA���	$~�>�C7dP�hj���?��a�������=i@���^U�>��Q��E��₈����i-M�P6}<���P�4Qj�~ATSQ>��p'D��J�u��U���>	P$�U]ۇjzک[p�9�$J �n��N�D��2��,#��tzƈ ���ӖW��ET$����%��	�5t�JQ��>���u����r����.&��J�v��l��F%<�*��.���<Ra��&8e��؏Q;�H�2v�S��|Vs�����O���޻{��6}M����υ��"��_�A�&�2���O�ݡ��Q�,~˘mD�!m��P=��,��`=��7�ɴC�aۏ��I�,�=�-�E�hZ9�5*�Իν��p?4��|\���?vxv�٤����H�ʉ�2�	�Y�ma��5 Y�$�~��ݩx�j_���{M��m+<n��l�B!Ө��J I�Qb��y�3Ѭ�e����xP6�ꄽ��
R�$ּCVi�<)�=����)�G�<�E$�^y����]L��bz0$u��D���%�r,��i{Qwpb[�x��w�B�%T�puR��rF%�!0�J�u���R@�覱v����M����^�D�?9�2p����2���W=�i5�5n}/�<~m�`)���%��̀�e�~Z��p˒��o4�Y^���_K���v[��.+ T����6�y�E������'�ޡr��T���2�����J���W7�w�b��4����!�cԆ�%�/�R�^b$�LM_�u�7�B�P�ѻr:�`mTl�-�xn���]46\�@B�q��X���f%M����q�cs�Vgh�
��qΈ�gr�s̳��/��pΙ;Յ�M��pKp��
��p>��̏����.	���C��Wb����3=�B��0 �;�F	̓�㽁|V�ϻ��&>V�d���a`�.����s�JȐ}YOQX�v���SvPn�z��O�����8��v�F�t(��}�kun�A��Z�� �_X��R4f�(�M&�y��V�ߘ^b��L��̢м4p-?����Ly�iϚ�,�b]�$�c&p��i�����W ���&�/�|D�rT�T9h��Ϳ��3�����![��z7�h#&Y���B��0;�L0��c��q�SZ(Y��(�e�'Kd�˝�ȝ�b���[C�Q�_�6��Nm�銯��+���z��Et�����B��ltD�P�-r!FSԖ�O�Аuq}tE�?V�����v���a6Z��B�%�%�ŗ���f4wk�C-�'����:�G�PA8���k��(J�_`9$n0���׺�8u�u�l���)?�O��b0,���}Kx3{s�ᘺ�"�X��b�����"����Ym��o�h�}�t�H>p[�ʽ�e�y��F�'��h���׼~���a�'Zwn��g)���p��������7n{
8�,)+�"NM�~��Y�O>�HIe`��|�LCf��dk|�6�D���Vd�p�2TQG�u�4h�b���?!��	
V#��HJ�&��!LsDvH���a��C��u��o(�Zd��J����bh������K+�,��ךۊ��]�	V�]BN��C�|%�l�-�D�1)v1�����<"�D��>��r*�H�M�E��;�J�!��iU
<�X����B�5�|��i� #��Ou��L��9/v$d�u����_z���B��mW�%xU-��ճ���,�G�_��D�o������y��J�̙�p���N�_8N���L�Pj{X���*B��)�o�>4S�xE��$���g�Hi.5�<�	�Nj�5ٲ4.+��þ��Ɓ�NjG���Vʶa�'Ue	>�Mvy#ۻ������r�����n�xk��E%E"ye�BtY��m�eZUpkE�����ӭ�W��jՆ�ȓ��U�z�#����T����̃�C��4��)�����j�Rt쌉Čc�a�ZH������Y�ŵܰ�As�������P��I�xYGhIT#��vP�� �`-F�"�ti��2��}Ome��Sx4�5J����o8�J?�º=��.�kZ�0/-�Q�,Xd/�O�])|l��f�۬7�3�0����td�k���dE=�r���	�%%Y����Ҥ�W�Q��ès�(��~ ���8�����	�U+k ��Z	��_#qSWpD��*P3j����Q�r�IwƵ���n-���H���	��kQ��
����F�S�$�HJaLP兂��d��vh2d���\��� wl�������WN����r��qYC^��z�?�0��楧SƋA�Q%D�qϳ��x�$��;����
��g9���.�D��W���Ý��&�ҿr,�)���~�����H�g�XV$}����"���`�K2+!몁?�dx�S2TXiC!�TN$AEWC�Uj8���Y�����fTr���~�x��/�dR��]��U 2�p����f��ї�3$�N4��>J`�&���'	ӕ��ŏn�$*�$f��j!�Bvx0&m�+�};�2���]��WY�mKX�rߗw%��_%��rB���V��_�e��z?�^A����tމi�������Q�#Dh!*�Y�W��7>��+�049�(b)�k �AZ��E�ɻZF�	M[�Ȕ����U���?	M��\�4�E��e8P/�78�h�+C�:�uRs=;��Nl��B��Ѧ��+eIy�E#Q�:7X�dtL9!�h#e�#��m��)�V��_�W\v�lXŚ�fB��)	�)���	lMf�)3d����jM��c
qA�!�ف�[)������e'��C���q�/QU#�ՠ���x։t���]��(d`�	�l��E��=�[ �ᄪJ--�B����S��xv+!�.p�n@�7$�@�:�W5������KBd�x%��<���/v�*�-�E��J���f蔒�nQ/=tRCI��ҍ��  a �� o@�����[���Z��:g�}Μ�����y�R�f�˾�M#��ih���l4 NEhY�~ ��s�S�NYV���}�5�}����[	[P�_��A����t��^:D㇘��h�g[�?P� eG�f��3#�7����BǞ �q�&�[�p��ŉ`eK��3�l�?�7҃��V���E=RJ��0n��rYh�
��/�Ԣ1n��B��߫9eMOY���b�;bƺ�HxH��I�@��HpɅ$u��7��`����'c&�ߚ:��1�>��7�9�W��S�덑�:�8��[��օ��lΚ,~C�og�tj�WdC��Lb�#sĩ�`N��{�o�v,�Ѵ��'�+aw���x����&R�g�$A�7��Y�2�^rG����A�>$��[��\2tp� ��(aA�W��V����̧x��"��)߭���mȜ�=��LĆ:m�L�/]��+Go6r8�=q�l���G(�����F
B�+sޏ|��d�z�����W�UM���&���`���J6eӼY���ZN���X�_���&����.�sN�]lXF�9~�������_��F�.��̩�p?aN;-R!��v�rSxm��1�⩽��BI����w�6r�B�*��[�������1����$`�F�7l���4�v�ܳ)A�3���>�G�ꩱ�NR��k?\�eY�3)��F+:�뢚�>��Aސb�:���Gc�U��l�V��'��Vx��1| ���v����`����]`��,>�������ȩa��!B%��(.!��?��%��-�s�vbN��͛$(yJA��0sX�so^,���h�A��Ќ�S2|�c,fW��ߐ�w'�#J4[���ۤ+�n]��(�4[��Ol���Q�g*�l���O���FӖ3�)m��B�lNJ�'��X��[�<�9E)��H�c����4��p�Ԡ��_�is�T
��(�T��|��#)�֬7{�]�Q~E|�'g�rl�`� �8%_�O�����ipp]F���v^lF�|W�����"|n@�u~��M���y�ޝ��%8J��ѻ��z�w�c�㮦�e8�(4�������\�e���ZM���)�����:#%�4��/�䤇��Q�T�{��X���������3o����Js�+�G[�g�AcM�)�2n8|���]��Ds����u�}j�aX��%>Eȭ$�ϦCG*�s�~x�dsO�ҿJ�u�,�ʠ#ۡ��lb����d�*Z���������:�ȝA�=�ԙgR��$�9pm_��R�zi!iq���i���2��Z�:��&�wBg������/��t��)D;���'ސ�N�Z$�eI�p�4��7lV�����Op���8�C'P|�%������q�Tq�'}Gfk��� �j�0�c@��{�{�0h\��o.���2!����+��EMٕ�`��;B;\����?�U�i�dg�u��y��9��"F��G�Pk�[%'`;��=���H%�o��_ά����e��3��g��37Cۋdq(ϝX�eľ�ȕ��?m����1=�P�"'T�k�="�� x���^��8a��o^�1�k�i����B���Tu8�� N�C|���U1ٓh�Gϳ�|��̃\E�aN���<k}#�p&���*oϫ>>��ОѺ�1���43y�6R3y	����R	��&�o0��Oa��J���L��RU�V?�n�&q�\1ݻ$F�rgB�m7�*��` �N)�&H�ɸ�/B�/t[QZ��˩�+^6� {�~F))�Rit���8�����1�C�]"5��x]�;����#`��8d� ;@�����G\`��[��e����۶�8~ j>�t�`V�0�ٴ���;�k{��<W���%�\��tDڹn��M�}Crȓ�e]6��EHx;�ױ����w�	e'"�z��Y�8���O�$�ML�B���;��;�}2���p��AՏ�r�eJ�t���uA��C�c��9�/�Vy�J����<��+E@���B5V�Uus�Y���Cia?�cmc����i���)e��O1��&�m^�SBh�<U�6dyC�c�Xg�g-ەH����?UY�8x� �c4���i�ّ��u��(fB�L�ܹ^4�z9�[�f�:�_j���p�V��$a���n��A��U��?i�ei����r�%S�����^%>Ƃ*�o��X�b" �qZ��?�Nf-�D~AV�o4<7i�7��q945\[Q2<��5��}��m�ؘ9 o����2<cNUUB{��l5�Y�X/��E"�P� ��ޠmYҐ8�"���j�cb�c,��uj���?�@�<AÒg�b9n�m��f��ײ*´��oΈ�[q{����k�U=��M����3Eq��,�F��\slQ�� ^@�k�L�k�7O��4У�Ώ��̓��ޠJ�ӂ�2S�.���rd�|�֖�a��?�����RM�[��H[6������R}��Jrh�KҘɊ��=��E��c�_�`�/MjQev��X;e�o��X7���]ZK=���xG��H
1b�-�t&Ec&�-晖�g�����}�x�ދ�.�&"�9���S�s��r�:���J4ʣ��	��/��F�J�p�\nH/^����>��N���+Uu��e�à�Ԥ6��Fs�s��t��4g^*|����:0��NgB��2_�}F ��K��%�#�U��N����8�FKR����U��f��+���J���O����;��6=����T��_��]2�GI�aGU�j���kVK�"����N������&
߿;ֽ�w�b�kGn.�9�"�����>�o�<E��&��Ey��:�lwH�@:�e͗
�Z�����Et`z7vڻ������b1��s�U��g�R�{����A�d�����T�M�׮=]���9{�a�6ø�n)rK}�4'�[u���t�"O��0,;�0�Tt�ŵUf�*ig��3xi�����D,��˪��8�0�P��?��_qwZ����>Ұh���eo�O�-w��i��  ��"���G�u��:����	*="�c��DA*`�Sָ��O�l��}�ڡk�/��M��Z�u(k��7 E�nܸ�2=��=��%Y�,�����'���L����_Ȣ� ���9�4���&f};�eYx�sK�e3�y���S�V�|�yX�aDbZ,W�&����f���~Н��i�Sz����oBC�_eD�R��.��;A  �1j�<�KnS��E��l��տ-�.~�H�TBK�G�Ϟ�	
��ܳ&~��x�G�?�������]��r�W�ò�����F�v)�
� �1u�Qi6v�T�&���>�ګ���V��o@�vD�+J\���5��������������<L�"Ů�+� �d83QM	yV΢�k?<������)�����˯�1��ͰAyj@��r����v�Hĉ�⭚Yx^5Ez�1����l+Y{�s����Ů���*����#PA-px�:S�5�g�?,
������U�r�KKEv�j�g�}�;����Ld=µM���e�d�3���&�M�����`7�7���Q��S�]�gb�_�����ޟ`���C���L�ט��Ϙ��J��Y�!̢4L���7,�K��5:�㟛��.�WD�3��T_)�?x��i8��Y�C��ԯNIL�������%����^A���=�e,\�>��v\m�cPx���Tq�wϝG���Ӻa"����u;��J��x��V�h��n.v8\O>�J]
����̌Ie&�wg�kV�D �U�NR����N2^j���G�5r2�'��E�ZM;���\�m�ZD�Zc�������{"�_��~��'U�����n�e] Y�+d~��V�����E�7���nS�ʜG̢X���s�ͬ*�j�^
D�A�$���������̏���Qփ���}�){�Y��N���Ε�v��@��0���4g���v��}���Z��(q1t��"�E�'��Zӣ�\�HZS�G\�B���n��Q����<��}h�PS)f�^��p�b�dgR���nS�"ID����s�0�Z���g�;�#�9��̼/c��*�v�M�e'�x�U�jǚE���3�O?t�@-3a��KY�M��l}[�7g
�����?U<�sI*��%��@���O v���ݤ� ��Y�d�Dc���sB��_b����?�K�"���6ƍ4���e#��P�ě��Z8�b�1%|+���%�`�@�:��.#���1F�1־Wp�M�4�x%%�1���M�;�SǴ>�XlS߲���x��q���[b�4�;rN!7?�J�]P"�M�_�X����?݇k���l�Ao��JK�"?P׼�����I`\�7�Q�7�{b0h[�4$��U�6MzQ��c�d�>�a�$�X��2�����l����A�N�,�	�]n��Ю0����j6v��P�a��)A���Y����I��1\T�EUj:��mZ�-	Ud�=a~Tq�̽Sԗ�Q��Rx�U��1�upv����MA���lB(���G3FT�#n��W�""Ù;�Pf���q��v�#Z���s?'b���9�|7�ȉ��vJaY ��y���S�u)�\����0��B��p�,��}.��&/��lV�̽"z>�i����̛�%�aֆ�����w�i�O1T����|]%��
PL`\�t��m!-�L�L��M��L#�bu�;��S��W(i�y��:_�Ŏ����@F%��e�<U]����"��LtF:�5���iyL䴕��{}�*'���ި=ך0Ň���IrBP����u��^��0w����W�I�>9�������Y1F�cTM�Q(vJ�/O�f�����3�W�=ѥ�6樉��s���N�2������X���A�Re���[g2���>��}�Qb�4x��[��$�4�C�[&�2��I5m�~?ƾ�s��;�/xA�	?���?����s� �i��	)8(8[�oY��F*d���=�&8S�<��0E]j0�)�E�uC��4����x|���4�+�`�n��A����Rg~�>�c,\8�	g�UI���?�j��>�<a~:Ҋn)�I���E�o�?ܯ{�-��Y)�1�4��t}���ƌ#�*���_ FF��R��v���^"��sܴ�Lޚ�(qK\&�W�u���X����^�C�	���RFS�6w��"�pzYN��7��ŊDqXgvS�B)K-�bf���(ӽF(C̈" ɑ#w��j��V�Z�B��!�<c#��x�+n}�^���$>?��Y�m���N� D*uW��\�����ri\ۼۀ,(ҧ@�Fk�p�)(�s��V��p��i�����fҰm._��&|�^��w'}��F�x�4�ANA�,��Q�3Ԇ�h2�������b��'!L��m���rRM�~��)�y5 :P	�vq;�a��a&/�N���!��ئP6��D���_ūvPq�wy�ލ� N6�ᦒ��I8���dx�ӣ����!ɦbESi�g�+M�!�庂� x��1h�N	���R\+��F�������&z��&�q1�U<&q�XY�7k&zM4ֆg�+jb��#mkl W��x2%����P�.���l�����DC>��~�:" G���[ku ��n�����d�MÑ�/D@���Y犘uoѹ�6�`��i��H�k�94���p��D�� �٠-KR�
�F_�gb�FBI ZpO��������PɋS�%�{���� �!��^
/t�	"_��O	�\x��E�n�����m�|��R�zս��#ӯ��>@�_"b���ު�z�`��j�64o�Fh�����h��OO{�<jZ*'���iu;�ɼJ"G�
o�N�ɀN���	�}��c=Y�O����	V��E۝x4����yÓ�[�n�8B�`��������y�:�A�!p}��?(.��7�����އu
����m�R�"lǔ��4�d`LWً��}�qT�(>���,2��L����R�K5ՠ�A�
\ҿ@Z�H��BI��2$<k�����DNl�4� �򀢙�?�6vUQ�\��WY�D����?�@�����T	�Rx��X�����F��t���������yk�W�����Dcm�MF�fZdE��bI����op�d���u�f��a��{+l�*�C�3z
�f�J��tc]�>c�oZ�.(�
�;�E��PA�J�L��繟�э(y`��-K*1���`�(��ʨ�%!xd�mA���I��`*�Á��+�^큏�P�(_��
�g�޹����E~�6�;fo�����b��]i�a�A܀�&���Ȼ9S���_��Ӑi[��ɷ�ְe1XSg�r|�?�tNx�f�m����KUIG6�Q[�9�G���k�s,NN�)����E�o�/(.����C���%�Dʩ./6��?zL��|�'��.d�.Bm���l�z'�Z��*)�TV��L�#�p�U�6gmt�¿Е��%jb���q���>��J/Ufn#�^n�t-E���^�d$%�f�	���Z<Dg�f]�*���$J���,�+�>�=��1����Y�{���F9>���o9q)��R�~?��x)UW��~��I�R��	��_.4L���&n$���R,DÛ�j�����z��Ԝ#�iLf��w���q:
���R��i�a
���#Æ��������[�j
x����%����:��nG�a�7��3��4���i%ξXFҲ��@⭇;�?3�c]�|�鐔�+�Ջm���.�{#�,W�]�'��ǉU�هM��z��_e���}۴�L���f��)�-i9c��m�u��\��蜽&y/|���<������a�C�ڢ�����R:�<�*�q�zy_�!��\<O��;�������I���g��ȯ��ߣ#�I��=��H6�n���ӳ"��p��]4���p�Y��@��cd��Hwe^�?��o����V��ihC@��:.�$t�Y�o�?
l�/[K��w��?m��Cl5᳕ά�k����B��0fB�S���������A�}ͯEyhСC���u{I`����3.��Ģ1=d�_䠠�Z�ƹ�/X������H=l�=�ģ���J�2P����9DI�����0��R�فvi!�S�oF�.NI��N2s3�K�Q�p�B���fN��Κp��!�v�z�,k'�\�O�Al�+s�[1l��V�_��a�Q� կ�����n�cm{�	u)Q�H'.���H���@VHl��F�5�����;"��[y����Y�CIo�5�Z�ҍMp�����6U�f �����g:� 4����E��i�y�5��P�3�)����3��
�0���ǮhtEM�\���c��n�.7��;�T�`��@���_�(����l@��ʂ{��m+H`���/q�]ٺZIa�Y /ܟ�%�� �S0��[2����R|B{&?�^��^��VR�����$��Qt1_�]f�����fUp��ԝ���H�"�%T�)# �?F��:�7�W�Z����F+�i�H��Z6Δ͍����V�Ŭ�8��
/�sH:9.��h|-YZa:!|�\dIJ��K?�hP���*���"�������R�M?��ś�VѦ	�p�^itm�v�&T?̙fap8�CBW����*3B�������l�q� m3��1n�bb��k;�F�XW2ː�1���}q��ޚdFw'9�Ü��*�R������F��UtS���.���eD%a씘)F!�р�+�+��eb��D���Wz�]��y��o�q��E�V�W���am����﹐�_�/�o G�3�nP��'�ε~N��t�<C�Ћ�S{Y�sk�Q.|P�E��F�$\`����^�G7]aԮ'?W�}��dd�̇�1�[�#����$���æW~�w;r�����T�Ұ��\0?F�-kJ��I[Y����&�l�E$��OCE^��3������o�Ͼ��)< �m�_)�J���*s�4U�!{��H&ϱ�7)�Π�6�v=Y$�m�7��&>Y'���e�l?<#�@.�,@�z�]�D@�?�iI<Q��E�1��&^�R{�/4���.��|�<�R^5��))�2�j0��.o8g�>2�j�2���A�l%�K`��y�w)�j�q��T�q���aq)6�ǅ��Y�����d�cS�I��oF��O���A�
�Vut8[�t�Mw2�z��g ZQZ��ݐ���s�0D�+Vs�#�G���7��ݔ�P~�V{	�uta�`|�U�1n��Gf��0O�f�dQ��&�ö�.ɫf7��w�2*\��ns�|+C!�<�����&]zB�Hvɞ�'D�EW���\$�)%mg����� >œ�Ei�o�_��4S����3���_�_��O��;r;��@�ЩN�K;pR���0������L����Ǟ<R��"`rs}w;g���B�Z�82N����%�^L����撎d����X����Udy�Gu�S)E��)�
4�.�?n���VN�;��5H�B�p$y��	�J	!FŸŗ��7`�0���	ϭ�=+w�=���O��������.[d!�?�6���'1�p��=����
urhd�h�L������x��l�s7.�em-��e���4ʰK�Ne�}O�r@�
Oٜ^P�+D���P�l�G��gH;8�b�|��@$�Q��ta��Y˥+
&>P�y��]J/�O���n��d�٨J��C�V|�`�F��k���Sp������`�f�t,̅(����kbf�CA��Fr>o�{rР8iP���V77h�]�W9$ �j^KL�~����~G��e��dr����*;b�锯6���^�3R~DE{DE(=���A����D*lDCw����O���'\�g�x%�L���#�����'0��f�<�ߐ;c-����݀.�j1�]WХM��selö%��� �O�.��;��+�;�p��Օ,�>��P��:�[����¥��/k�&���>��"��ښ����X��.�ȗ���OG�G>�P��;s9i�
r����V��%���`�V-[@���.K���m�
��u��Bi�)^Ƚ�̫d�ô�W�(������'#�ҏpR��{%b���%�i�X�W��p��bd#@�-��D+�0����2����O��G:�g_�^��Aǫ�?g�6� =b�H��'Z�� �Af$�H4�\Q�Z��
���(�R���7g��2��G#?�]�68ݼ;i�d��%��USJ�j����3�<�B���,kO�ފ`�93�fq,�L=�n*P}�8G�sYkc�l�-C�x��>�*W�G]�H���`�ָ4o����\�$�"L��@]���K��(���� \�Ȥ��R:g����1��#M�Q�f��9�۱����N��*��ݖ+�q�Z�'��B�(��fx���y��Z�Q�1粙�%{�����R;��D;6�F��H�l$��>�����i̒Fj�K��d0<�I˫� ���L1�eVJ���㈫�wn�H2�T���;˘*��k�p#ijIK)z\��'7y��;Ͼ~�~DS8��Y��g �Sս������oR�#~7/��n�K8�sOO5�ڭ5���,��lN�b�e6���vw�L;��<�bt*�E�>N�w�f�JؐF�1V!W{F
��'=�^8��s����2�hCkM�t��^�g�"a9��z0��_4ć.�á1��(b)�"�������t�
37���ٰ�����ɻ?�w���Ҥ&y�9#���+(J`X�RVn7h�dX�LI�{�a�s��L��J�����[L(���!9@J;�:�H�ek�N6��z3������w�ma>Gң�A���]�n ��p%gÅdس�H�>ʦ�OA�Vd|2����W�t6�����d��!�?S|׹�b��ޒe1��T�k�V��9=2y���v:�� ���Z� ���D���d��ؕ�o��W��G ÷K�(ؓyQ�wG�i˔�����4v�)���P�p�0{���h(��j�����B�C��&����5 �OϚ��VX���ȃ����n�T�����%xm��S;Ե�7}s#�o� ��x�??'<��v�~��KUuG62Q[�7rF������hDΗR-���f�wv>��ž�VFI�P�;��^�F�C�����؎)��󢒩N�RF��]�����o3�����#٩��6t� �^�|�zԞpM�^ʳ+��Q��x�2��w-0,��3x��Ak������ ��y��{��k�W���<�$�]��U�kp�䱒��u�ю�!�N��N�qTos�S)�K|��y��f �m�%��ߋ��ZL��I�Q�Y��p�q!��
6���=J�U2��+����K���|d|�[}3W6�H
�K�C�m3��RlX���H�����w�2QuB<e��F0��n��נ�=�4i��Q�VO��P]�镹�"�㍞����l�s�w �8��	���%׮�䉛v'{PLXb�mR�u������Ga;q��
��_��Yfx'��)�uA�	u��F&$��H�fW������6����w��4�Z��d� ����Q�奱��l"��#��"}��zz���~��L������٧��`��BK;r�Ԟu5���J˲������nӳ|s'�����*��Jv'�69�[�U�X~��Ͽ����x�6Gsv�N����F�ף�:ɢ֨뉣'D9)Jv�hXP�HN�_n��n��A�`t��Ӷt'g9���0������F�EY+�1��ˋ7�x�S'[J�a=��.Q�s�4_�˦��}?ϱ��f^��+���v	����+O�̥ؔ�g��b�(6�����}-��ux��`h|՗���y�a VV�xg�Q"e��A��n������~{�2��>����? �~Q�5z�I��`�~�L��@��d=|r��d��`���W�5�޾O�6���q�O��a������kD�����_L�|ѓ�}_���I����:�"|$zgC�u��1V�_&�=T$��� [�k^���|��^���Z���t��Ǌ�����D�,��$��� ��a؅3(\E�/
T���4<�w����4z���zJ�[ �o��]ޑ��s�����I����[���ȓ��}����ϙ�Q�Nx�u=�B�2Q3���_�P&�d����!��1���G'F��2��^����$�<X�Z�&0f�����ߟ*wM؟��P���*��r�~	�(r��k����_�>Ə�"�ޞ�^m�������G���ST�'b��i���Q��A.�Z,�h{m�����N#����o���vZ�6���F	��)��g�X�O
B�bt�h�L��ʏ��6K��
��I���/��#��]�&�I/�oVd����ؿ��B���v�K�����ZJav���'�~�3�d���0^õ����O�G���>�^$�h�.�q��mq����Y��ٲ��l�[�ӷ��!w��t��fu�򖧐/ϙ�~`�M|9�I�s�L���nj���҈e믯c�I&��r����ǈn��_�`�,o�>G�����Y�lU�aѾ��Lfd��4_9�ZY��1n��,��+��Ӆ��w�92�v8]K����ǥ��%Ӈ���J���*-JF>�)n���=OI��U��wz��#��,_}'t��s|���R!�k<��+�)���_�q��ړd�oH�O�
����u1�T��gUL�\X���tj��2y�����w<Xկ>lK��u0��H�"s�O�A�l��.j��a�Q�V���̰�k�=h��;۪�z���޻qS5��Q����j������''�!O��!)���Q>Ĝ$ f��Q��k��|'��-�w��@���7��|�zk�A익���������G��E���$��y�-�Ϲ�"|=�����V�G���;��z��>V�e�x������+�xV��e��y�E�
Q�Hm�ň��X4�ӬY�;oW��U��.�QE~gŗ��?ocDBnR�{*o���ό���$k���%��L��o��7���nō��R\y"�󕝒ރJ���U!uG=��c(�"�S9��P���g�wL���J��@E��aF���>ʏ�r�I�p���r��kd.8ٖ�k���/�"<J�6\]��{0m��"F�9�+܊ՙ��Z�p��-̪�:n��_�	JTa��])Y-O��O*ħ�)�{Iw<�ao[�k�x�#������9���SFs�f\Ot���l��,�	�f���l�W��&Z%s5i�k��ɊOՐ��M�&E.h�X>IQ�9Q�I;4���0�w�d�_�z�����t%��9KgG������(�"PJ.-6�t�%<3kۡ�m��/�iK-E���!��g}�O�	�����9��h�T���	<�;i{��}%���ޡp^�V#k#·�hsR�Ʊ��9��=�)�3�9-�X�h
+���=��B�g���n�x��n.��px������L`�����3��*���>�G���8��uQ����M4�V����u��yl��Ν|�0�sdB� �����W����e�vHג������|�t���T[_��A�x��z"�$I�g�شY�d˴2s7 cwG��S��1c��a9�3���c/�Fv��kʄn�}J����0+-��i�{�x����C�LU�-����"�2��H,�+ND��3�
~'��l�&O!O#%�x���g]�|����e�t��;�Rx��Z˅��[�y��f[��*إ��d�/Z�.7Z4 8"��$cZ�r2�v]R�M̓>l"g��_�}�z3Fdک���/s����]<��~J��\��e�RQ9����D��sdTD^Y�*�z���h�[�x���v�u�uYWf��X� W�	��=Fzg!�NF�É�a)�ue�U�t�o!�P��i��Uh�e�ڗ�8��c87�8O4�#~��)�ؼo a���J�5���U�wُ�����G���
L��JY�l2����bSN���
!N��r���r��!q�5&k���c��x��X}��X��^�
d�Go4Ky��(*�����.����v���$k'�o
�t|)�z�������Ǐ�QqW��`�B�,�%	�S�q�-չ��~7ŷPY���"�!����/X��Z�#9����v�Uz�֜2�B�9�E=��o��^oy��m�g�U��U#��+/~ҥ?��'9l�:�ɰv����9��u�A�(�l�pя��nġ^�U������:��ĸl~�'Ψ���D:(��g��Ncj�Z-уdX%�9c1�MĨM�B$���z��
�LU�� n����7�Ƀ�麺�X�K��jf�#�`��۴8�~�_�o���ɣ ����;�T�#KSoY+�X\mTI'殽xSM�M��윆�̂�\b���L^^��ZtRW�QY( �����b���e���)}�T��*�)J�V�0���Z�J����|%�W�q��a�����E��ǃ��I*���,>^���7=�J���>X��/9|M*>�h��({Qy?G
����^m�Q����^�>�`^�U�kD:�up|�W_l���Р	 K�;�����=g0��Uu��ݑ0�U���t��J�nF��xI}�d��y(��d$�`��]���2�{�9�|b�u͉��|g�H��b�b[�+qF�~SrQ��OEo�����?gwet�&_���>����Q�oȶ�O%��4}��_Z�9Ɗ|Ҿ;va ��H۝�&Xy���{*��,�c,�!��ɡ�[���#6���۷�կ��
���w�D��"�iC���-��ѝ�"��ⷷ(A9�H��� ��i�s�	���ی�KJ���
�?ޤ���E"rU�=­q�R�qK���m�������g���T9ة\BR�Q�z/�����އ�vW�M� ׉����]F�m
��K)5�6�ʶ���-s�T�pqEZ=�Z��%�IQ㛫� ͽ�*$ޫ�`�� Dd�&�ۊ�<�q��k�H����0��9+�9Ww�{H��x|�Gw�	��!�VB�{b����,t���NV��2b>�쬸�F�b�ea:u5��)P=�Q|��m�G
]���=���X�#<�KmK�����hاQ,�@�X��<�x�����*}\��������ڥ���l��d�@���a?��*<UB)�Ϭ�񃟼)j��ӗ$�#x�f���X�;�m��X�E�2>`�֢�������-��e�~�����R��/�ט�6�D:k��)YT�M�Ss޲�6kG��g��Z��؈YY"���:����+�X�q�G�Wae���E��3����n5TՇ���/x�0�ÕM��AD�!�h�u@�M�Ǎ��ƨ�����B�@���@�Nh1�����y�o��3��¬9����j�^��Y:���(��18oc.;�Z�TTl�ʕ�v�d�1��]A�*X}M�7r��s�.�A��@ǋ���+�v'_���z@��A�dr����睖��@d_B��À�7Yk�ֈ�cϚঀ6z�&O�K�������G��t�����3cJ9QW��騤:��r�-�����8������q��~���#��Z���m~����Z��l�asI�O�~�B/ELZ���f���f&roj^=���&���_����]��������� /;��,��c������D��%����Vt,ѫ#4l��)W^��:�Q��hDb7����4�gej?z�^[-��d����`Z�7n��s���� 明OEQWh�K.ͤ�Pz�f��_<~�e��&�=��MTӼ:���`H�9�
4��s~��KT�0�y�L�k�����lĽӑ���p�Ё�ϕ�x�M�T�{�c��E�)�üm8څ�ǟ��l�=�fEt�^b��/R��!.N��o�=�SUZ�%��إ6`�n&��[G۝ŋ���ɴ��}��['k��T�����%���H�Wȹ�w7�$6�v0s�Gv�%F�q	:ʎ�$�o����tw�FF45y7谮�\��t��!/��T����Zi��W��I��A�R���x"w-n�4�4
�����,��VsiK>2���M�Q���8rC����ݸ���T�Ƚt���!xZN��{�dc���gyz_%�iM�jU
�(/�iut����]p��W����4�D��XW[N�wb:��ks��e}�m�\��}`��~c���x�63��^8�)T�z��x(%9C �M������E�8��Rw/b$F�-EM[^O��a&P1���!|�5D3_w���[#n��H���������>��Gx~���08��C�`�j������B�-B�B�!%���I�9��fgl��E�8i#�\y��;�U������n�P��TX��ճ�u��� �>䷵(���y:��yq�u����|{�ŽY�����oĲ�*Ի����|��i�GU��zt!�ߥ�c�{�
#��O��w�Y�q���w���:�aP��� w?x�/q:M�|7��W9/��dV��)v��<�(j[�|���\�ToS���i7#s�<����0���;��	���c��a���w�3�T�c7j^�4O�I�韠���9�~ۧy��u�ؑ��D.]6����[s�6���{���ӛ�u������f�n-
:GQi��<R�E6����>��ɲ'�M�'P��Vw�.�ۦ�����cތ
]s�xP�>ۉ���B�P�����;Bl�R�{*�矊�L�HSI���됋�f��u�3تzq�3l�����ۋ���Vj��T>Xd���C	�R%*����MMb�z?N�7����,����W&dZ��`=nvWJ����n��Z#�(r�&{Z�x<f5��2jW���s�w�=�z��vӬ��`����+��7!���o;�Om\F�T 7���XR�e�4<�P�x��;�/1w<Hs�^���R]CV��2?ʨ�a�Ŋ+SD��8����>�G~��}��9E�����6u���LۢwFA���8�x2�gO1
;��
�!`/�w�5�L�3�-�KvD,ay���>5t��ʽ|]Ј���ހ`x�*�6������x�5^׋�w�k\-]�C���j�ʇ'��U�x_C-Т\���p��l�%���$�Q�����'Y\�5���x	t��W��[�!����553�_�~
��n�#�"�J��g�l����KynV�<l�v(*���P��C��Ƀ��Ń��؟�)�Tߝ�0�q� �܈ �['��	f�:ڤ�=���u�����H�BE
3��h%c0O~H�N�\���M%����p\N�����)�*R�<��*IԖ�W�A�ۺ������՗���˽~˛*�i�haps˄�*Y<��Ϟ�p�~�������9�y���Lna���g?|��5`0k�d�Ҍ��?9��h59[MZ[�>_�F��ϡ��v5q�BU%;���"��)G<�M����njD}�m؞��+�vK�{��f1�ʊ�#E�g/[Z=�v��\��n�\J0y��xV���iEP��|���n|a\�H�e��(��A%�B�p?�gOJ_���f�M	��B���mٚ�"�wڻ��>B6�m��=�q�ّ��KӚ�����4�hF�V&=�Mx���b$�b�8�5�M���'2-d92}�e*� Td���px�U|������YF����J�Q�3�JN�i�V0��H���������f�c����KXgSE�y.�8F�"FH{��hO�����$���߬����"���S��i������J�B���|��!��<Wg��1K+� ��"�PM��FH�*�vs� ����t*�r��J�̶�CBlwoF�nئ�"V�K�R�������|`_X��R[���Z�\p͗b~i�j��%��G$Py�U��!� T �{M�Y.��֑��h����'�.j��W�C:F5i/)���_R#�ѭ+��_Y]|�A���%{�<�v�^p#���O�P"�i�cp�5��K�!3ƒT�`j�q~-FN�,��a��a�ژͷ��:�?��y�� ���?�f��TM�6[g��5��^���Q7��	�XI@�1�B������;ӻUmx>5a.b����b�f���?�w˨���m�qwwwwwwww'��@pw��Npi��-x�{B� A��侟�]�Y3g���}����]�w]�޻�	{Q��ͳ�<wmù�!�/�}�W�	A4���l艿 �x����B=��%������-G���m�C�֚�鎯|�P؀	a9z�$y�>�,ҡ5��`,�;��y,���>�wM��n�
�0v�7��E�[�M��d�a����.4j�����d�07H2[��`�����A���m�ݞ�if�Y�z������g 2c����7A{�.�JR��p��R�S��f�Al���F�+��� n%�9�XׇϷ-��k7��|-��� �v7�n�xI�VJ��3��l��o<�<�ib���UW��)��tp�A���afۭ����U�i׸j�e��c|O��Q0Oh��xH�/˺!hf�a}���8�/ÈI��$l~瀅f�SjF�Y� �)�S�2���?�@����DBN���%�(��=��-�
��/��q�-�*�  ���
*�����BN���ǎ�xc�}��@��
� �'��Z�z����-X�9b����B�+v��>��A�塥7U�<����л�����k��Rp����.�9���B�˽}k�Ay7{7
������B���M�[-t~�!��~��h5��JU��hv�k_c�����"�v��V�Fv/�V>��å�TF�V���X�JW��ow��S�s
�9m������}���ˈ���t��p$p��.�m�7�Ã��P���p:_!��˽�M䭤�S�8�9��"�7� ^�Sr����m�k4�5�Y��\ٙ��W�	��:�3�� G���:��W�.�ҵ`?鿡p"%��)`+�i��¤���DF���W0� �ȑR�ivw�Ex7���cY�J��W�,�㵭�I
��|��ԱSI̝���Co,��j���'��wH<zG���XW�ƞ���|���Jɒ��������"���A��J�C�Թ����x6P��O�2��F�_��(���py�Q��s�������U�.�Rb�>`c���ӟ��_Z[�Z;���wR��JS�~764��6B��D�A�qE4RR��&�w�P�WO���)$[¦Ow��>�wЖ�6�����4��G^�ܘ��ؙ�Y��N�k����DM"����'�*�����әJȃ!�d̈́����L��h&50<�P�x�f�)A��w�@Y��(�okiK�3�boS��/����b�&�\E���Vc���\�U�4IQ�i�}|癆�;���%)�R�/�@����Zv���U���t�S��v��o�~V�Ρ?��A�����֟x��`l���� ��.��|�����P��� �$����Ɵ��'��KSэ㵲�5��^!5��d���ׅ8(N��~u��Y%��u�)@MAx�`���45�CǤgVQD=�ZCc�^�=��_}��X�+��V�π;S��@�su�v	[aݰA��z��LNi�FZ�44^>�����c��(��1J�!�˟ۏOF5���Z��(��T�0���N��h���k~q�E��l�s9��a>�T+�`%5.p�y)�;���7���J�nR�a[�r�ՌV�
K?��԰���Bva�1�����xe�A<�=$A�|�b8%<�,��^օ�]�J�߬�E�@�(C9Ml�`2�øa�L���C���4�9�Ee�!9�I�l�f|��)H��H�UF�M�5���q$9n� i=���\þ�����-<0N/ӓ�5X7�����<�� k� #q�Z��v����[~hr�m�-��*���H�6�+O�+���b���m����1<&�s�W*��ۓ�(B(X��Ԓ��o��=��2���=4r�Ĥ��?�4�}D�|Gp�!}�3�w�&�o�͟X� P�2��6��-�&�8dbĺ��@��[h�Q��F���2&�U���� �斂v�}	�$K��?p��ǘ�b��;�lyB���^����M׮<@sW<��z�����D��ۼ#�~���J&q�����1	�'��:+)*'���eu�H�a�w:�����O���zb��9L'��s5˙{�ZG�&�U����s0̹=��X�t��6+�Kd���e�*|�済�$�������z�
;��U��-��zwIA<�iĝ���,�t����P�m;[��S��5�$h���:�A%X|�+���M�K˨8n�0�������aX1���,��|md�O���	�G�<��OX]��g{-�h�Y�D��V�1����%p�Yh�����������WP�'%���_?OM�* ��wvM��М�����Q�T�<5P̈����m=���A֊Q1�-(]��}�61�^��+R{�F�onb ��ߨ�U����?��F�ݽ�9�q�C��Q��$<t���Ð���Q�����$1�Z䶶���yɯN(����qr�(��	H�h?�)2��lX��v���k/���
<˺&�N<kq���s�h�ᎱH�t	{��,��+9�N����Ȧa�BR��˒\9>\��NX�mA�A$�ni�bXd<r�Ӏ�U���3�
lk�4��{!��,��Q�&������ƀ��D�.o壯��y��a�V%� �g�vY��?H�t9�#W���9ϊʚ���9����&]��Fk�b�D�dM\I*�G�O�Q����c1P�)#�A㹵K�V���v�D��"f���'�Fz*{<�K���M4���6��Kv��rc��+����P74������f�C�z��i��9$�N���v?�K�C���]"�5��B���6�!���G�-����zO��M�e~�R!�57)(���~x#���/�F���ɦ���3A��v��L0�z������@8`S�RM�ß,)������oz�ɁV�HaF �,�ǍVQ��P�)}��Zy�􋏗ΰ��ȎBJzI��͑1������w2bٗ$u��hemAHi:*Å|��6j�	���B��K����c�h�k�����t_;}�(>o�8�ij��㬷;���/"�C#D�{Y���50�;)�/՞���1��Q�J��l�[ie�m�OZ�/����Qs��)H�
`�j�g�zs�MAE*������3Ҏ����yv�!V�[�f�;���[\i&j/�or���<Xr29�G&p�A4�o��z ��	K���>ￅ����".�CY�k�#��^�I�%�\��y�O� ���Y��K}���!��������]<p�Ff��a���RW��W��l��E�CG_�SDj�]t�"F �ShgYarDtS�?[���R�,b�J���k�X��ߠ�]X�N�V[L�䂓m'�e�,a�����*�M�"�4k�(t�aڽ¦��L�����kbF�Z�>�����D�pɞ=`��SHx���s��l�`y�]�����z�����`&��(x�La���#/;f�׺wF�9�N�.���蚖�2�:�"��~ܬ��~�������/��l�UhkI�dɡ�u6��S4*��8�t�[�����j�iAz�ى �&�@�w1�!�^ ��߹s���^�f:�^-�8TWGS��O9��
~9��� 8{��P�eU[X��3��U���Ov���[ �K�%���]�H��{l��I̼�	�`"/�������I ^{�[vD�hɶ�p7Ͽ�R�I/��i\}8�S�'#��m���
�X+��YYS]��dPj!1�?�qk��Y��h���>�z6��$ԍ�<��]��C�k�$\���c�%��(���B\Ֆ�N��7���ձ^n~��3�4�k�G)��i��q�o�	Y�~TS�f�#
F�P��%f���«���\�5�}g2!��>�K�(�:>��]�J�Ƕ�
��������4TQ*P��#� 6�R`ׁ����G:�0_;tR*l��YE�d�+M9�	�K^�Ql�ˑ�=l��gY���os'�����վ�ȋ��J���
���'�L��l"G�m��XV��9��2bU�����#�\:]Z, #!Pr���AF�ir�O��gӫ���&�!���gevz��>~-��BAo�r��W�lafa��2�"t����aw:=���W�`�f�Z�N����Z�l-��%,(<|k���{��Z���]�3��MU���\�������M�󯗮e������������|n�t�ژ���`"<x��~Y\#E>%x#����#�:#����ܗ+���~�ң30�?�j�s��%~��9sH�qo��y�g@�
1CUS99|��S�
�RR��cT�!6o���@�♴�鐓���6�芾�S��aC��v'���S׻���(�"�$-�?��=��z��4�~����i��CNL��S�eR{!������3�{�x�π5�����7�/b��%!6Gȟ�0po%:�n1��X�m�3�?p���a�p�
���h�f�R�3�rroP|��\�����QM��)7%�i��d�B ���?X��Y��p"��E��3���Z}��,����h?�E��;�����:*U���/胝Z�U_nZO�3X����!��PW�	�{���ץ���|�Z.����_vT��\�����]tW:@
�x�ğ�9���n�����e�qﯯ�;;M�7��v}�j~�C�����H��:+���P�礸9+�|��d�8�~sv*%������+vJ�W���33C�l}5?��,�u��'}&x�֫��+:��� A��P?���91�d9���-.�������g@���SWLK �Ϫqe������6����p\۬��I����e�Ѹ��l��c�Oھ��?OZ�{� fC+7t��?�C�c�{��.�&_�%5F@��=�R�����k���P���ѣ�����ê� ��~�9�$�O՟>�axz��U��y'�)�"�e��ժK�QI�I̽.Z1��?_�|r�ap'�qg|���S����~q�%������v�st��62�e�^/��|7�pі��;�7R�Kx�
Ư;ݨ�0�Eo[��9� �9��1n�ƸT�b+�����h_K���6��=��46�0&Q�r[d��e��#A��C��9�M\7���[85�a�w�fe����uT�n(	f3�����[_`�����,\�y��R�=�g���̦���ۑ{@��pI�/�S�,Fy^	��ZFW�O��������m�,|�_�ѾP��M�h�@�������8�|Sc�s�ɒ��'���w�ML�B���1ϺܕŻ��j�O���N#=�;�0��z����d;C3�l]|ټ�T(�Ͽ!|`A�bޘ6����h��Lf+>3.>Re��z�;}ջ� �g #Zp�p|.��Q����|�����ȺGP=�,���F��!m(����8�oY�{]�Q���Q|�Cgr2���^C��w1�wi c�|�ep��O��6h)Rk3&N��uF�"�-Z�sG��!� G�Vg_������4�s���!~���sˇ|�O��Уg����>R��XN�B1�s�Kcru�,駭[:�w�pr���ˋ�D"�<a��Z�`����Ƌ|\[���K�.�?7��L\}"��*2΁�ѷ�x���>�GSnn�2/[y4�ҦG�ǃW)�:��b�2�����k�� �t�#��;�[F���Z�he������ȐQ5�4"F\v8R��Z�?���M�H�B]y�w�����i� q��6V�$q���?5������Ai�Ό�������"Z��e�=���Z8���IE���G�嘞�D��5��;"G��tP� ]OK�5��A1O�#�s����Fɷ��-#MM>C%g#�t��h=�H���o� ���b7lKF�|n�P���O��"Ia�,���@oJ��e�\�=Vς��^7|��59��00�b���~�I��޺3�!?fA�y�;��XЩ��ޢ����F����vm��>��?����W�AQ���as���k����'7^��姑��q~
U�*^M�����z�S��P�?�
�����~�{��!�B��V��Ň���ۭ� *  	����uQ��J�VH*�f�z�z&��dڰ�����9�X�ΎeB���:w�zPZ8��6�}��r3���]g�
Ӟ.�����3<��6��2�i��>�w#� �b���la���CKIW��7J�{_26��V�����ئe=چ˷�g�t���2��H�}7 ������S;�Fp���^�����oB���`ހ�Ԍ�k��+Ԍ9ui�I�dpyJ��%cL�x�{�b�_oЁ�+�qjDz敵�ڷ{n�[���6�i���l5�%s�y
��^��w6g %�ɰ
;?\@�E�W�Z�ti������<4b)���XV�����b+��K�]�z�.b1 ~Aԓv�*-/ru�F�T���}V�DI��y��pV���Ո^p|�g������� Flp����4}��ܘ;9���a3�2��I�2�i�zԍ�H��4��&M��̟�g�q�di��A��`d��|�d:֖gX�L�����f���Ę�|v��ً�Jɯ�����3���	6�^�����geRIo����(�\�S��l����bQ1� ��0&:H�q���y�i�q�K	X�%ܦ0c|�W�]n��)�����QH��+�ѕ��#"\�C�k�s�bYq[lɎ`Ŗ���n�PͿTS��O���/��8�r��A���?���I��f*ҹ�x��n$���Pw�S�v�h�e���	���i�i�[��&EY��e�w���¨5�����V %�b��:),�e��2yO�\ن}ȣx�W��3��%ý�NZ�'[ũg �g50m2��,�=��֢QT*�!W"2��(���ňo�������=a�G5}�����"8�\�����m���?E�p��Y9Gͻ5(Y�w:��C;�i�#�qċ�6ʞ�	U�R��j��O�	2�ݙU�BY9w��q��4�	�X������_#��*���_]��8	�6�o�IKh�.(��
H�H>��Z���)���cj�3�$��5�9܁�UMON,B����e,��v-_h� ���]~s�P�
�sC�I�Xfk��v��0���KV�����u��C�����/�8�{���E匮g��Tvg:���}#�@�HP"��9�sb��K��p>Ӊ[d�.�:a"EB�p�~��-����.�
uI�
���w)���D<U�
��E�k��UV�"�%ޯ�o�� �Bv}�|�9�H��ov/wopk��͈J�IXon�Rqݏ�U_"礪P�����a��k�rH]�}�(��+��_Xޕ`���;�hY&3�pӲ�t�.?V���Wǉ z��?85��8�GR�3�#ܙ��'S1��a9�8�Or麏��.�.q`�3{P_Kwe`��䈊�]�@�:�'G���@��|L@q������ ������� +��X�Zp��������1PN�p4��`�F�Ydw��P7\�C�K��B�D��6M����[�9�j������� rI�~��ʋ
��4�a�c�<�"Y[��/�Ϫ*f��!��'a�;�ػ��}�̈́�N�.���s	[������ۡ�!�Sr9���2M~I���Y�t���o�22X]��E�^��iB��	>�f%�}�"3��fb�`�};u�(�<�e���	0�У����F6�Ò7}:�����Q�r2f&`"ۜ={2������+�Ƭ�ic�7s�oϾ=�])މꆻp>�a����@E�������Z/l��-Ս��K�]�+�Y`�,.�ǴGR%�Y�R���A�>�6.c++�\��� .��F���f8Y�l~�`��P�Y^��g@1��uӘ��
jT]���٧�Cly��CՃ6Nm�0*üH8�z������*��E����`|r8%0�d���'����X/�uM��4�_D��L��q��0��g!Mמ�M�/J�ޓ���/���ؖ�p�i�k`A�'aUX�T���[C����
5}+
 �"S���HAY���Q%�((�^z�4\�h����T�O���	Nz��lGL�C���� ��6���`�U��fS�Ş�I���j�g�Z"0]�I�*0��0+{�4`�H���}Y�)UM��;���{u{�㽎������/V{������,0�	����f��,�Z��g����5���`S���Z�h��G6��[_��-��%�3�P����!tPk=�|Z�y$��,��Py�ik��mQ��Yˏ_�X��X�an�rf��X��%z��5���K��Z�+�e���w�����bzH����/�����T/�h�K��O%.1��~��[�6�t�lF�Ԙ�s뙲^xDx�Ba����cG�m�N6��f���$�NJR�H�3�|4�h��o�/T�t�2�Ŭu_~e:'�c-�yV��ʊ�r�e�Ǌ���[�4;�X�ѯ.h����e�l�vS��2<2s��ds2����p�ү)K��i|�:F��U^��!%֌'����7��n���W��G�� �a�~���3��P�@��ߩTLt�.��*�/\�p�X���dqA/���Ax��lе�R�A��ۘNmL�.u��Gde�
��,]8vr��o��:�x
V��u���d��h�ٷYsAHI5��W E��8��ۘ(�T>���oMDxb�z�r�G�5���KD��m��l�W7Y�l���!enge[��B�{�������.&�S��~3��j�T��V[˼�]�o^�I0%t�'�7oV�M��n����j��$��$���1Du&[Ʀܲq����$��2��1���B�^{���!�C�����D$�x_�y	I�0��]�:i� '��(�_K,Pfy���WÀ�����Bi�����8!�ᓡ����uz���]�~���h쐿����Xί�Z�0�M���J!u���/�@c��#�!�nƙ�K'Wٱ#&�L%�q�OLA�c�+>
?F�)_x'�y�_v���wm<u J���9#A��M��Oa��ĭdG��Dh]�%����e��X�`�Vxf|�u;����2f��2lw}'����B���M����(9�����q�������:(n����+�KU����l�
�r��s>�$��i<�M��$QI]�����M�y���8��h1:����R)�X^�b��L%�[��g�U�ev�t��_�8Y�4�B6׌	Oˑ�ңx�	J��2BQ1��J~�ءov	�ԽZͲg��lPM���9B�B�����`�C��~�=ɛ���줿�:K�s�c�ȴ������؅�W�X��)�(R�$1��\�js���UV���é│Qu��Q}����#�G�C�!�?;�Sj�02���F6s$$'g^��V�G&1��Mo����У{���!F����1,����5�F[�)�t�y�E����.ځ�A��CM�o�xЍ"�7��pY�߇�0�gq���A.�<6<,�9�|k4+"��OD�wj��7g���ң�F�t.dH9e]}����{�3��跣��h��Ɓ�>'Xb ������|������/%��4�iSsA-���z#��?�I5XMPOh|�C�[����6��� �)LU���ݼ/�}Qh��:,�������m���ǁ���X��@�#��yRJ%��l{�E6��N�a;"H�NdC���rN��6��ޙ� 5�
��ȥ��$+z�wcDȬ�Y'���y�������4�Hx��1!�:J9�\\�P �;F��ѝ@��2�i꡼?j�M�ꁞrM��Hϗ�T�|�U�^7k���������3.�+Ќ���=�i��h���L��	��T�����n�	�M��O��o��N>��̶��LD����H`�q��	��u�ԟ�MP�g�?�������ӓ/��~�O�{Cz60=�a��-?�s����	3��8�C�۹E��گ;���
��|�_�&�l��7�!|��i��VM��2�'��,����Nz{�
�,�~?B]����N�{t��-Dw@�A�K��3�mk�Ug����/��;
��n�"�  ���1���'s��oh��I���_�;��̙}��p(���Y=W���Wmfs``A�d��?ЖU���
�F�ii�%�:����ˢ���FEoުL���F�ײ�&�u"X��n���U'+���� ����K3  �֬T�a�d#l�e�WagI�zt]����͜���Д\�d�&��Lu�Qɍ��GU��[����]��ƀa�s��D���q�ۘs.�gF�J�?�qr) rO��1'F��ĥ�`A�h X5./��?p쑁|�e�[���e<a<�����m�M��M���l�{��,}7ٟ�A� ���o�/��s�$�S�f	��`���c����M&������]iei�X��\��^���1F�j�n#If����M��PLoT:����F1�����i�sH���=I�k\�6UIQ�vIl��[O~���,ȃßEh��Z&�.H�pc�����M���MC'ʈ�zG}p�nW\�O0#��00��@J����(��n��Bh�[1A��n��B�[D}��y�~�G�����,πws��"Sr�HV���v�!���� �ط�/�Ǧ2���_�(�Fe�8�v�P�윪�m9��9ժ6iN"{���*ѥ��Sg~�Ԧ�O�����_��b���(��S�]�f��yáҏv�+���o������s<�P��{*�<�6Z��Sޯ��5O� �{�A41N�nx_�X�D��:�`�br�?fL��M:?�!u}�q�)���g�O%θ/�D�88�[�U�E�h�(��'�~n~��lo5pm-rc���������b��� ��B�qٷ��6��tv,s\�
O�J�Q��oWZ7���bhL��Rt�٢�,��z\$UԄ �0T��OJăy5R��p9�1��K<D� �c]mr�4����͛}z�c��Q�����yЇ2��T/��~�CW�Ӏ��qs8�4ΕB�����Ó�/�"�����BrҠt��A��m�Oq��j�}��zK���A��W�!�� ���+ݥ�j�!l��U�ܴ���xi`$S-+8s���)$0�_2�����󩺢�"����U"e~|G���ti�θ�u��-�F1� ��F:$hk��!.Zq�>_���׹�������?E�����e���}��L ����~����i/<���  �@��j�3��?�썢�p-�~�n��>L�����r���M,hk��8M�s���4�[�}���/v\|�n�K�v%�!W0��/�J�=�6�#�
�z=0E��N⫞�m��l ��<~�e�=����[��uy��7&���) ��;u��~�3�YdMH�yb�,����mM���Z����$��=3c��	_�E�B��l�`����C�K�NՑl|��R'���2OJ��|��_����s����i,�#�:`���Q�VI~���/mE~�~z��U�d3�;e�m�Ȍp��� ǩ9*^l��ԃ�,�H�r\�Rw�J�uv�-RӰ^�&6��"bP(ҝ�*i6�D?�^f�z*��E�V+�N��F�b5���t��I49�8^ͳ&��?��ֶzJB�(p�>����Q]�e��.�S:��41��>�����=�x��pG.E��m	�o��(O쪈�C�@PW:W�+��2R64 �@O�����L�ԖL[�Y�iy
�����u{�z��GN�t>{\J����)Fs,��<*��@��D� L1_`{יB�EJ' �N㓷�9��e���o3�nq��!�D�Ւ�	��;��Mփ���.����}�1��=<�չ3s/)
��ԎH�;�R�X���߈`�\��b�����<��LR<�ʺ"��o�Bo�/��@�[���h�k�_�R���<�ά��D�Y{�M����RB8����	s�H����w���ad,��f���� �Q2!~�@���1�p�Kz�r�FeA�"�6qx��MN~�r}�n���s�yد/�U@֑�v��L,��4����Oo͖�p�X��3�j�sEn�R32i�Ӣ�Hje�X�k-�,o�Hܗ���Y���=qNDP�r�RW`<+X7>�l��e�����	�̎�v�A�BwU� ���ȅ��6�{s�$��y�E�l��a`J�o~�&�<�%%a�K�V����q�LW���5����?��W,��,��0�n���y�;T�_��֋.�C�D'�;B4*Q���:���=�;�M�5�jE*������V��v����:��x�ʷ���ϸ�$��ڶ��G<>#�W�R��6����~�N�Z�d���_l��7��Ί����?����^7�Y��{4��C�/�v`��="x��d��\�g&w�J<��i�Z�M�lAby�����χ$���	{�L����c!�H�?M�p�S�C�l
��Ea*��`S$3Q67m&0��\���_
^0C��B�d�뻘������ǅ�����v:ι�ߧ�� k�R>��#��n|��>X!��Ɛ��ɣA�?���V�����#�W��Vz��2�^��(�yEw�1S^�"�!L��䈂�X����x�Ž�_%�!��c��^m�^2�(�BxA��[�n	]����b��W�>S��	4Hm"��L{�T$�II��x��V��	�5�4���&�lMF�V���Ҝ�%#����j��)�P�V�Tc��Up=��
U�s�&(����+��biWyV՛�� ^k�F���h֢x�N��o�qD�܏��M�+N�����x5Q����V�ȋ_̫8z>25�&�V�-M���7΁��꧜b� |�Q����Tw�"0E��dm4jn��g��xQ����;۪V��!v��:��|��IR���ճ����/w��&R� :�M$���>F��
μaLXAÁ`��t%�T�gF� b�=��� O7$I�C�K�|�K9��5�q�X���D��B�b���dwv���.�m*�G��&�B�I����%LQ�ޞ'���v�1�e]����պpK��]#*@F�P�qV\&W��&�Zg_��q�p�D�7���g0[o>|��ق0�h�K��B���+�ҋ�Ǜ�}�)�#R�zޙ#tCI����ԡ��T^�^��g�����+�iХ�������@�m��������+�m��]� *��?8[����B�46\�5h4�8KXC��7��IN2�uN��8��\f%������N0ijTt?4�:�!�=XQʔ8�����soe�����Y7��@K�2��ʜq�L?AbF^�َ�y+NU�<P��<DG@E�~PT=Y�S���g��nB����˯6�a��e�r�ڊPv����%w�<���nۋ�5<ͥ^͇|�^�n�Wrh�[/�ݖX:��tc�3�$��d����_R�I�3����2%�G�K�[V<�i����8' ����~@�cV���Y�Nu6L�}2׬��ʌ����������{Q��qn��g��םJ��5�S���2��Ye���
��9���쉯�V�ʜ����	a�;�����?]#P(��7쮛�`9�����|Zܣ�㊾�^0}C/J����9��(�>(|n	�x��{�䔶* L�^��ئ��GYn@"���)o{����|��5���~�{��z ���n����j��`�r>����vo��`�#ٛ8�z'����kED��Q:.��yeچ��+�v%h ֽ�@�\4<���j����癑���~��w�����m���D�2���:�6�(��L�Y�Eu����WE�᜿��%N�	R�k��[�e>lg[�!y�(����'�A"򠐦<Ä��v���ݜyHէy��l\�/�ǖ�ke����F��8�EGg���nUQ�r�em����]�V%�o����0�j	ʹ��=rA�pR	�ۤ`��3�;"'�9���O,�jԄ���T���Q��1�O�4B8r��TW�ht�=Q��}�"(e�6���m���l�
��K���)fk�ш$31;�����nmIfsν�1	t@�l�zjyG��x��o���Ǯd��
^"��h�1l-,��t���~$xq���2����%��� �����܏i@�b�F� �����Ob�������xW#.ҟ�>�an[Ϯ<��{M�ߕNec�e�a�p�a Z����x|ܐ[d9fg�_{���2�\���D_��*9>��9�8��d?��>M�Hؾ2�@��)����8��+��6��^@���z��v���v8�z�'qǗ=K��<�{z�����ԜbL�u~���%�iO�T	C;,0�n�ڤ�^���$5�ʍ=����hxhh2�ɆW�^d�1�9��]EX8���΋z�-�ˡ[���I�M��=�NhJ���*zX%9@��s�����(:��!t�1ǏVbB��nܠ�g��2O��.�
�,l*�'��� >^�A�4�p9Cʆp](�>T��ky.4(ꒉ�P���s��/�4�n>�dX,�/�4���u������DF?=�퀄����!� dw/�j,_T��*�'�+U��қ��RZ��%���73�)`%mS�#����e�Ց�S'=�rR�!^��k]��:��|�ѕ�Ph̄m6����f�\yy�������`�W��uט�4a�k���닣 �L���T�e@�V��RKG�fK���t�	�4�0��i�5Ǳ��$tu3���0�4J[��oXަ�
�e�؎k���^}�`ƙ,q&|�D�B�\Y���@�,�u�S�,�j)��y�m\ś�]kJ �?�m(_��n׃�[���)�f��v���v6�g�쇀B���%_����0|>�L��z�w����横(c+.\�����Ӧ*�2Ո�J�hف�g	U<g�w�T�Ϳ<:�O&#:�d�,���.>H#���8k���_������L���g��7�tA�X#���~&�1%�o�[�z2����G`t,0y��������)<L"�9�ջ�)���h!K�G��pa�5�|2U�Y��cPk��������*�d@�ձhk�UY���cz��r��q0�@(�����kq]�v��O~��s��(��� ����X�q��i<wz]�h_]y�X�cpO3�k�5'��g.���F�C������y?8�����r����*�y���Y;G��\�������j"
.R4ޏ4���!�#��eu��	�*�55�e�X���P����2!AS��?N^<���eO�@d�M�%�.W�J��W�(��N���	xVM�%t���)%��o f����C��|�fF�Q�iB�k-q�M9��ڱD�$�8��9C�MH��S�#�_rv/�]Z�[�����vNX�X.�8�<�쨽3\hH���˥i!��A�GWT���ƽ'�[=ڋh�t� NLN��H��Z�sPDE��{tP�1 � 3@E٥�ߢW�����D��k:�mq��¾Gc^.�.UC��R�_Yͯ���	���qR�.S���g�>+�����|�p��E&���4P0Or�[#�?eḧ́�a�; �M,q����p��2�v�2�d(�7�$s'����c����f���V�����@�s�2�#dȆ�H��us7���6��=P�����!XV�"���Ωӿ.G��ٱ�]�3�3@�v�vǒc"��!}YQA �?Ma�{J$H��!�Q@lZfI�Ae��m��Μ��d�ѥ���vP���eP�s����9�Y�g)v˒6�a�-�R|���c�lM�y�P@�1������bl>��'D�^c�	x�B���U
�K�Ῑ�?����JN���3`�#kg�zL�����b��v�8v�"���/��n��n�*�T�#�����ѐT�i`��\�<����I�a7�ࡒ�\{#�.&r�����;ӑp�~���YU8�H�2p�棽����kJ6�s�A'��0�$��i�#�㧣��1�m��<��xni��m�)�1�;�9d�ɜ�s��r�U&����h��G)�(�(G�W!�,T�Tvk'��"�2�fq�	��+l������ӷ���"d�ٝU+��F�J2V�o)\ApђCr5�g��n�PErs��ÓA�����W�lw~��MsD��^�*���h�nU�L���K���zT����Z� �l��V�f�\��}�q-3�#j"/��-ɗ�G��e>�G�F
�]�,��zE�Eْ���A��~�"�aD��YB�4��"�#�\���bD5�%�^	2>ʕ���T�U8ٌ<-���5���4��C���"tc���������A�������2o�u׼!���#��zᔚUT���*�o1�?��i�����FC�xU�z�n_5��6v	�V�Z���� cG�bS�`��� ��/�bG-+ϩ��!��u.��1���6ԉ�(ZDU�ڑ.w�ޘ�7�t=�}̟���Sl`��{Y�P�Sx�ft���c�%�㹓%����Y�3�����}	�N���F��*LV�t����P\�ݝ�RE��� � �墙}�kT=���g�Mf�w��%
3i�jS�JENY�7k}��)��!I��U'AT#��7���Ǫ:Y��oo/����AVȮ!F����H`v�Z�/0|�����h<K�<��pm��k��Ma��"v�%������̥0!��KjrP�$x�!z��W�h���ts]QMm�:��ޫ���C�^�H'G�z3R	H�`@ H�"U�"�bhҤ���T�ß ϸ��}�/w�1�v�Xsf���Y���P�F[W���2�ǔ^�Z���\
�p�.�M�W�Pt#tc���oJs
H�h�~��_4/���d�$ጦd�{��U��Q�;Ls�kȭ�r�TD��+ݐ�xQ��*7�	U���Y�7{~7� ~�kW!����o��F�����	�X������_�\�wGI!=+�DbSV�z���	n�qv�Ȍ^�8C���{0�m$t����US�Ϭ�@���]�V��s.n�)=����(DM`�B����r���圏�?l�Wx?V��P1Ԉy�#3\|��J��W%yln���뱫9tJ_K��Qyc��ܣ�V��Z�[��z�HV����_П��"4�x2W:$�,��L�g�k�?��bec�΍̌�'��)'�]�5�6ޟ:�<@��\�A��'���r�
�<Nn~�Q��=���dM���X���8=ʨ���Hb�PzXU�d�/���m��a�%𫔘�c�VD\����L+�������1�����	\�����yx62J��Jw��O%�&u�1Tr;HCQj?`����D�@�:�S�h�:������Š�r�+w���1n���:'��i[�����aNJ�*�������ɞ�4>�����v�H��O��-�]F��df.a���U�bl:��x�Gߙd%�s��\&JΆ����Ц��)�X�@��'���\�1J��ХX9��mp(�W�0��Q� �i1�(���%kY�ύ��������b�Z�`��
<X���=�ʮ�h����71��ϰ1���}�{B�}��[b&]~`���Z�Me�����Ҽ�B_X����T����\_��u�0�n���|�s
��/����g��~����L�x�%�v�ZW�%a6����� �iW��U����Y����vX󥒚�A���'��m���k���7��/z�I�,�eݺ��'�#`��-��u(�Cv�4�d죉�+���,�z7�T����#�L>$��@
�9\�q�M���Mkߊ��jwY�|A��Qq�T��,f��s�H��Q�d_�Un.WϦ�3���ͫ������7TL����{ʾ���xE3<�+DY~9�%�DYp*��L���0��T���Adxs�9�e�G3��������
�m䲬^)�-ʆ��BZXU��]&T�K��!����;��5�F�q��SX"Yֱ�$����~�k���D���Hz�M��&+�nN�Z��)
��~V�m3����,Ӯ8)M�{�@�X�JZ��1�/�ʰ���8�������wՅzW��q����u��1&�J^�2xPqX��{��� ���D5��}��_Ĵ�6A����Z�
u)�[rJhA�5��N�n�s�.��ԉ�c�c� e��}��|�� [�t��P->ͼ1��Aw���I|�n�K����qJ����B�t}5z�&R9�y���/B�NIA� �8M�e��]}E}��u�1��R=�G���"�M�w��'�(�#�sOoT>��_���4d5�9ړT�ǚT������>=�����v�:�����Gđ&��`׸	۾9��Y�,`��]�2F�ݺ��S@Ž����y��) �')�{�=�A�9�� ��bL�0)�|�-��SzO�@���S ����Ŧ�����kǵ�,/pN@�L�GN��>_(�U��
ql�KP:�^:i��'@�D�hg��:$�yk�ME�p|f���CzzB7���M�2%`�Ԣ�#)���O\���Y6�j��,�P���	Bl�3�q]�=#PIj��d�h��ƹ>�����'�?�dlsv?�����ĸ���e8�j�b��<w��UDE�6�9!��x��Q&��eg>+ �N9��wc�ዳ7�f�D����]]��G��ô���`�W��}Ñ��Z�ޱ�^N�Yd<�Ĭ-a�{�(�
�^�/1AeŨ�lx�]���H���1+|�O�������'5$W������nk����a��K*l����.�Vŕ�Sr}+X�{�	�Ͷ���4<�Q}Z�x�8!K#��S0���܅f��c�H��zJ�
OF����������>��/�%Wt=�Ό��.��+&�ܲ4��Q2ҫf���`�j�ϻ3]���'P�;=b���D��ķ��U�Q�f�����t�<���.��[�F{��r����>�4�� ��u�>R뗃�/�:x��>�A|<��S�*'�a����Y2�v]6�$���cJ�\Ѹ`ѷl/���]��q��:���-�+}��տF���T;� ��]j�yc��~<3^�c\ÉrP�J���Y_�f�*b)��?�M�8	&ｓdZ�Ԏ�����/�T�$co2�ʌ<�m-�f>��\��]qJ���*f��&b<}J��㬷����ˎt����__T<۠�U��*�NT=� TʞC�ޓn��l!�*��y�GOYd�x��xݺ!q~蛫�R��=���Ia�̒����l#�ΔDj��fLXr�����,���n�'+���G�|���ؚ�z6I!�H ��K��V�fS�h�- �ӉCf�\�ޢ��vyO^����ٴJqyerq�N����͉�9�%�����_�2����%[��'f�y��A�Cm�.����[T�����Z&8�	K��	N�|y��6�W] O�3���1�H�|��?5I3�v=***�t?!�]��������&���ϛ�0\ک{[�b���X*(�ڦ*h岛��w�0k���S%�� vl-�#DB��_�41�텉��$���3���K_l^��6���%��h�ϫqֻ�^>fG��KV�_���"TuT,B�N�]�K7/`�.u}(T��m/l�qo��^ o�.��`��^g�) x��B^�?_�Wp�>��s(����[�Ǟ�Qc�p�C�E����V�}:�*��&�%���y]1t#�j�*,�:J=dS���b>0�:i�/����i2�!L� t�3���#�N�T�z_�Bz�y�ʎ�������mG�=���f��B��fk�kjǵ1��}���3���u���UZwq7���.���.#Q�С)��x�o�f&p� �@���F�HL�d9�څ�������)�u
 ~�jA`* ��ջ�zp?Hݢ�����n���(׻į>��Ҥ��E����z��Gk��ydy�k�1��3;V7{�����/+I�� ���7��h��>7/�r�
(�휥�L�bcc�<��aa���}$��s�����u���	Z��6��tVoF-y�1���xw$�g��V�����K��&���ד�dޞI{d�`��x8�G��3��'��-z�!�|����,��W�
�y�*�Q�����5������*���
]^6�����!~� =�D���u�$�u���CpP�)��v9�����j��Z}�����YJ1�H�Y��m��W(1� n��S@H��P�ޚNǷ4�EV�8\�l�~~Op$��]6��ܸ�lS�Zt��R�(��d�V���E}�����.*_�;z�I�)���ӱ���u��P�ym�P��_�����t��@�)�lI���o������k�R"h�, #�7yIu�`y��H������0�S���=g�Ȟ1�L?
V%����H��s���j�B��*����+g=��fo�������v��9[�K�ɾMG�����K��d�;���u�:������G�].������P @����4�Zt���4tf�i):���8`�C^��u�8���sN^����M�U��}-���͐���t��C��=HK�h��}n�3���pq�qU{��x���I��Q#�\����-|2N{��W�5A�)q���|�I��yC��I�Î"_�b��C�ly��ê���,i���ss����d��®��0.v���a��C�J�5���;�N*y� �ڕK*��Jv=�S �����o� ֟@�:�H`�{b�c��|����;>�D�^�^h��}�d���6&�y���g?pv>��j�8Z���Rw���­>��E��h��m�]������,�C}A�Uy0�1�р_ ��1x�г�lW[��F���A�]N-��+d���ޓ��w$�+n�*o��b�3;eBkU/\����"�������������/RU��X����;��ˮC���M�;ϥ?�F��*��Иn�:F~�	�K;{�*�Aq�b�W��j-�PL4iq�R�X*���C��ᮒP��<'O1�:[3�ϑ���B�ǅ}5W��AP���:��|����]��]� P�n*#7���p�F�`�)�(ؘ�	��1ơ��v����sP�"ȸ<T��ު��[0�+&|ӥ��Es�A�Ed�����}�qf��W��u#��|�y,iy}�ɪ��o�pR��%�E����i�'����9IY��P�_��ui2	���ߐ�۝(�w�O	�dR6���_�m=�t\��A�_kO�y-�R��<���֥>Dj7�1�R�d(�"0p�� ��S�:p�2�8c�|Q<�a#)�ެ�M�9xm��K2��Rnn�}u��
�n{�f�,�X,�)ML�p2�Itd�D��IW�$��;Bg����'s,Q�����'AJ��X�(�R�(��e����#Nm호�S��5���J�0"�n��5�9�F/���~�7�+��yG�gO#��[Q���6h��ݞ�>�~1X�	]?tD#��KK����Hk��������O￤e�4nl�,s0����ߥk�=��׀�0�������	gg��(z-Z����"&c���_f"��ݧ3�PK   �N�X����7  �  /   images/2b66d102-ef9e-4dde-8ee7-817842500f7b.png�XwPS��� R���PBU�!��B	M@E)R tH�J�^�JGH�.ҋ�PD�@QJ	
�}��͛�����:{�{�:���={�8c]����dddtp=��YD��
p6z�d�>��zh226�s���v�^"������dTg	�E2�3v����3 �)������7?�s��ܒ�G��/�?�مg��EAFv�o�{�/�}yU��..��=��} �����ɋ	�F��>/��-+�>�1�Z�%��|�����p%��9�#|*xPݎC��S<�'���o�9�^>�W1L�Q3����.�Q��Օ_||�*~d �֋��'uy��j.��9Z�*� �u��+�>E�� �U�L�.5!>�n���f��f�q�7Q�>��-g�_�T,�X_k����>�:�c;����F+��g?���r�q�1�����Uʰ���r�S[0'H0]l��?�הۖrm��O�������98��W�8
�}�)��;C��r��3���&��?�.���d��ƛ�d��M��X�2U:B�72���/l�b��!�#8����G��d�{��x���m������#럀�(����ū�e��}��� }�g�
�B�!��R�����R��QD��z�_/�)��1@�2���X�L�d �IQ�l���Fb� ��yg�W�o��t�Cy =�(/O2I)IGP�yYr����?"yd�{n�y�kΊI���;���!����jx{����QB�
�����8/�<$���9_�B{���H��w���;�a���S����!EK��ű���"���l�4kf�Z����Y�5h[Y���z�_Q59:�eɔ��5
�Iu��qV}��Ԕ��� ����TH��.���F���b�	�mM@&�cA��	�)�����mگ��wD��M]�_����Z�)"�P��R3���Õ�m��~�y� ���,[=lo��� ��8,�Lć5��63�*(L|�H�	�A8h-����"Ҍ*{D��e`ß�Cy ��g\.�PK���$CX���U����a0|�.Ȣo����G��EE���Ϟ1�$��|�B�ܵ[֘hkת���(k
E=��/��-,�$bb�MLc�虅�/�6R=xW��4����ZЋ'R�Uf�8n$Ⲷ���5]P�I1ِݰ�C�d��{I��M�7��B�!�P%�A�ml�A��ƀ��$�R�zi�pT$5h��h�p�V+d��<�~`pn�Ȋ����	@7=*谭��x8-	�v�'4k�߲t�]�Eo��ʍ���\~5c�U��-�Y�Ԅ ���D���҇ӌT�L�%�I<�X�(�,v����Wn��L4����P69����'8�r�rI(�d���`�G0�G�14�k�:���
��$(�;���lEo�y�B��^z. Ul����i��n?	���L�{���S�1'�:����\ϴj����^P".�� �]�@�d����|�� [l�T;���|^^�+}T�{Y=мJ��x��]V=�IS��7D������o{_le�@x�0<<�e�R
@��Ʀ��I�Z��W4'Vc{Jq�Ukg��ʀ=?%e0W�-�TT=�	�!�fy{o�-+#*�S�OH�)� k�F�,ѽ3�L}k���n���G_�,}^]�Ԉ{|������yο-*7����U�j~�afh\��^"��h�!�`؟�l��?�g�MMc�|�S���X{7�E��!�����r�~��ۜa_�}�p��&��D��%q:��~Wh���05����v�7��Qskk�
Qf㦡!�og�%�Β��V��t� ^�kp���v73�E$��F-v^�.�*r��NbX�z���>r��y�5���+�9���9�֫Ƣ�z�x��]�@��E�]���z=�N����%~�.��"h)+�ѿ���k�7�W�u�����e�⹠�1�}�?��V�v�@g�Y�a������%���כZ���a{?pt�n�3�j2\>�e(oí��8�*��e��CU�sf&�����3�R�o�^=���ǡ�^1Q:V�n�z'B]�4"Z�\5�zH\ݭ�1�q\7�2�H�}������������O������a�	k��\�1������ȷ'<��S��VئҵJ���`��lu�f���tAK�a*d�$����f����V�8�zK֓�z�V_C��kj�g�^�l�A0e7��F�e(�͝�ga�5��i��ʘWk��zT0�MH�	p�۴�f�Fƭ�EFF�W�4�z7�P2[��`st�c��:S�@C$R|z��X��#OG^%�/)�vr��i�	>�v0ʓ}��S�U�+�Nf��V?���[�M�RG�;�]��m�mG������2��;��pk-ǳM>`���`'��X��wTtB���X�g�/�+�4��Ȓҋg�c�Yh���.��7Q�0?���U�S�zw9W��C%�6�u�mƵb�0�+Y����������
H�h2����*u���Y�>(iS�(�ɷ����4B��u�Z+��0�����t)� � ]�I�	KoL
�l�y����)���L�whm��<��-��>��=z�$��"[#b'��9!��r�������OO�h��u��vuᑑ~_��i�����D�~CNS�z�흟J؍�Pfa�~�ϊ�xUk�2�K�� K�U5�B5t�F��z�ќ�l�zO���w.�{�oj��1�xlb>3��b��F�4˸�i�D���k7��UT�X6=Dv�O�Z�2��LJ�94, n��P���L �}���mu�����d�o�K ��p�s+�`�z�gup��,ڒ�J����o�)��6��u��dw6��m
�gf?���o���<M7(p,�b7�碨��_��נ��{�)�d��2y��z�ɛ�-�2�1�g�72�"�r����k/��g���hA6�.*����T��IA{�P�4|>i���7=�%^��0d����J՞+����y�:j�I�h8w�OT�n���^�^N�s|\CZ�劻�Kp�zY�3Q�):��źC݁
��ƌ 42ji�*�}S�!�"����0V-ӧ;��e���:k����U�d�w��[\ȯ��dzzz�>���e������ Ґ#	�Z��N>�����R:C������@����ki�����e���j��1�F��\���?�J�<Q{�rO�����B�1^'m�����A�d�X)9qc��ai�w�j�gN�隄�>s
�\����24������5:��(Ǌ���d-�ޓ�=���rT�,@,d��FU��E!:S~���5|c^�-;-���:���X�)�4�M���*�0J4��n��Pa��o���\��g��ե+�z�[�)�o����Aw�f�KpK3���蘏�<���Fi���O����3�ҝp����,`-V��͊�5���EQ�n���y�!Rey)�ҵ���վ��9��j��*��v���j�Ǒ�����`���=�&��h����8��-b6m<�I��nq��9��Zb��B%��[��n^��l�%�W�۶��O�����)���pa����M\̞A_ix�쑋 џ���^�!��&''g!��x���">�V/���1�__��-H>���`l�;!}0\��Ee}ˋ�n�y��:f˻�j�)��� x5�K����u�pu�F*;p����%�@p���Hj�W�Q\����W=��������X�����Uݒ���J����G��ٮ��J��� ���DB�ʾ�����4ܡ/���%$s��5�N�fj�m��$�_RYu-�*3�gdd�J��l܋�fz��ʪ[��'d�U5;��td�_��?��ų��i4���� /5~��&b�.e�"r��R�2�Ƅ�A��FE]��%2δ����7+�,)�<��N���։]�ϯ3"�u�R��y�<����h���g��A�hr�ʡ�A�W9(�&D&��7���L�Z��$Ξ�o%C)�`0Sg��L��m�g��u�`W�ISc��W�|Lc4?!�4�ֶ�R��$U-=�N����g�r]�B��pq�ʒ�32d((0��B �{�,l%N���F��s�Cw����_G��^ʰW���ǜ������tsSl��͖�ҹ�q��W_=�[�	F<���N�5�Fc#�A:�J��ҩ�%HP_O_����X�����Ș�[&����y�n�-A��C����6���w�(y����N�a[�<i6��w(��q���Ige� l�4n���I���V�Phfӎ��8�tw*)�����Mӯ]y��Ap���*���#�������4��bq���snE��u	\�V�i�/PK   �N�Xo�>��q  �q  /   images/2cd737db-51bc-41eb-8762-f3273c40eae5.png =@¿�PNG

   IHDR   d   �   J���   	pHYs  �X  �X{�M   tEXtSoftware ezgif.com�óX   5tEXtComment Converted with ezgif.com SVG to PNG converter,)�#  qIDATx���d�u�+wuu���9�LO�   $ DҴ��l�Ғ�//�����o˖,��%�f	H�� #@�<��9��t��s.�}^������*LWx�{O>��+�/�xF�`�5Ci��� ��ɂpE����0�(M� ~>�ؼ�Ϡ��E�h�slyh�lz�k�.����ޏa~?.�7*f$c躴W���8��F����kX'L�{�������������;��|O�ԏ�G��Iy�7�r��f�l�)��ϔ��_��R��zmU���˶ғgsy��YX�&ē�Af\|�j��,������XC�����B����c����
�k߅��,�๸zb$?wD|roS�r�$��%����׭�u���fHL��e>��0�w����q�W'3�����/��'�A�s&)+c1fL�0�y�����xP1�O�^j���-�^�^�1C�ɰ�q���K�pq�mȘ��r�H�z�Ɉ�3��e�:��U/��_R�|U�J��g?ٿT/a�}��=�^�׻�U��;��ں��>����Q8Jl�%���3����9�}`4
�JSN��蜼a&���~���� �qj5Rg𚚘�"dN���T���yo�x@�K�m��~u�fܱ��F�շ��jZj2��.M}�W̐{|���O�aځ��]?����m���w��+������돖s$f�݊P]����=����A�g䷅�Иn/1���V�O��߁�����͙MbN'(ok]g�V!.��%�7���PO99vje��M娭.��T&��&����1_XM��T&�Z�u7��²����Ȍ<��;]�/�^��_��n���y[gF��~��a��g�`�u,�!$��8��b��� �V3b���J�*��ho��4�W��^Ĥ'R ���4�Z�X�U�V�nW9��¸��]�82�dL��Ɂ2G	l6�.�z�Q��.��'W���D0���w�_B���������m��� oc�$�}B'�{��[�j��>���7�N����oe{�!(ťQ��/m�+a�P8_(
���:~9�O����5ÙV�հ�5msAL��KHnv�Q��t�l�� ��UR��1��.�t�Ӭt��V��`8F{U%&� CA_�41,c�g���/�h��"�X��AӮ���E���A%��"�_S>�&u8���ΐ{�k�z�q���i�����-�f�ɑIܮd�_�qkj]��d����"FYi)�������I��9,-�J�8�N�J&10�E8�+��E�(ä���9�X�xnIf�[�a�K����+aK�`���]�h/c:C��L[ZfDf|S�6/�.�������'S��T��<"Ay�����>̏#�b^¼���7C�PL##����`�8�ל�L)�a��d�d��yJV9�������p����_������H0Z�����[�������Zh4/�x�������TF�\r��p�e��lƺ:7�?�+�I=�'��=WE4����ai)�^�xj��e��D2�٫a��ӞP�?>'
��M,a8��A�#�Jǐ�]��8����A�uU��K����ك!�?�(�[��,8�+��8�N��[���Ħ�e�+�2��,��U�eQ�>y�,�͍5x��E�è0����@�W���U.~|c���*�Q���:�M�R^���"C2�)dm�I`6�5Q8��=~�vZ�J�a��#�?�}.4��3i��
Z� ��hi־>Z�E�9�ECi���9�F�/d�k!Ys1�a(� �l�P�L��T\-5�ƹ(��4*��̱83�3?���4e��$�:sB&�@ځ��2�sFe�L��,N�"ڮ�Z�I�.���nRք��8�a��	dсH%����Vem��]�z��M81<Y�3�$���i~���	���xlp>eyݿ���	*��u@�o-��S�#�P����U����ؤO�0���2Md�PVQU}7��~ e�b��Rq\<�.�~S��ȴs�V��*$��]��OO]Ƒ�qaC�5e�p�,�V�,�A3}�@>.ǂ�妭��ýsT�0S���3^�8�������Ճ7.�''/#O�t�.���!l�p#�l�[Mv-ҞLFP���>��z�S+�S�Ȑ�Qgv��(�6�:@���ذ�$�a\�tX�y��'����E�ꮀ�j��3.���|D�������[�aH����7:E� =�DzQ_��1b�9�ڱ�DF�X�8^�Ua��nU�e�HT_ ��U,c^�����(�����dZ9�a�[6���5X��~d2i���V�l��]"�↨�Dj��S�+�4�n�����_�4��f����m];p��	�	t�&#qE����كjFT�m����;wh��xbY��E��*Q_��\ex�^�>7�ya��S�6�`]W��w8J�?��/�]�82��2a��F	J���e���g�+��p5v�� d�zQ�әt��h�%�ؾ]�ӈP(�hTcHYY�_�hjߊ����zTK3����VR.�������.�(�b2��J��s�$��(�?��4�܍߹k��c��b������D�j��� ���h�C1�4Ӑ��(u�p$�Q�ʫܕ�(��Qj[V�y�Qf�b���Q�j���)T��g��t�θ���lu�ԘS�ȋJ0>�*�/.Y�7��ۡ��P�IV��h�L�+/E��G=�~�6��7�T�dX�7�Ջ,�3�7S�E�dõ05x��� >��M�EgS޹2�hքx&��o�����3�΀w!��t^���"��b|��G�P]ی��!�I�ӱX�hѼ�����_oǀ�����:3�ş������_|�nL�cP4-1��x��t2#J��,�d`��sIu�O���Y����2â�-��T0U�`^Q�~������?��K$k��2m�{��a�N7***�����0����d�R�f[���K��8~��X��.Tմ�>?.����e9��@M��><0����(�a������>�?P�Դ�U����R�5)�8}ދP$�&�҄��sJ6�d�(�:'�;�Y"J�_��:0��s�BPD}\Mʛ��ٿ��s�S��B�������h]w;*�u��o�^�Ao��Nq9�1r��I�<8{��ܝD<�DU\}G?$'�/}�&W9��=7(k"%v�����	���,�a�-�9J]��o�5s��S�B|#Ô�+�n�¿Ӵ�Nxb3��i�N���X<m ��/���_�f�_��d���2�_SVz���jS>�7��x83
�i8�er��X�#��I�Y9���4>@�/��0eՏ�,�h��\�_w�6��K���G�����sd����Y���T�[݁���3*O�xLZ)�ц������w�@\��i왨[����ʴ���B	��(5*�9Yۅ�����e�,t
9	��4�9)98��%��d����-x��i7FR�c���|{0ZQ�O�%��y^�d�Z��YA �U�m��o2%�H8Eg���=��Wˋ���-jA�F&٠��dm�|ҫ��Z+�rt��&��{�*%��)�t�?�s3j��sT�����R\q��.%Jq�P��;�2�GQdY+Sf,�1+�������VL��$�v����o߉py���rL�i�J����������[�8��r��|d�|�����&�n[638RjE|F����~�,���\/���%��>����)�rb!N&�^h����>Ҹa���>�jʚ�E��u�ߜ�~w3t�)6�s��
;��nI�&k�B+�[���s;�x��E�$G��\�tg�E�9�Xd�p�k�7�9�:sR�7c�xƦ���C9Y�<t�L��R��4�(TY�m�d�ErzlJnX����vqE�ߧM�¤��_
�CjcU��?��)�Z��F���9e8��I&����7"�Ί��O�4d���$�6%�ϔ����	�OŲ����+&q�ÏjG�� �Xg�6�$� OZ;�<V�0�̐��Ϣ���6��z�A˖�sX��\������|u�]��_��0'���qiZ��8��'��cq�"�L�T�����PT�}�����1�D-��XY�WN2N�jK���FG��r�:�co�/�k$<��MQ��ϸFqWMk�<��n1{#!�N����~|�ӆ��*rw[=�{�,.M������X��;�� �~�y�zK������oܲ����F����qyҏW����Y&��@����{v������僸��N��85�A��&"1��}�o�/���fū��3.{�V�����\3��V���h���^u��@5�4~��[��v�GQQ�CBJw�{������h�C��]� nq&��/���	���i��۾�D��79�暑)b~d�ZY��~�����=r'��{=~��ױ�wX�m�b8o��R~_�syXf�ya?��7I�W���1���{qcg~���xJ�<�$*����AyΕ�-��/Wҗn؈�/���=nSף�Ģ���ٖ3��W׿��Yy�!���,E�����:�АQ�����f�28��V�d�[8��p�)J��y��$ �ު��CD"��f�Z�vW���Vly
���Z%F1�XC1u��v�W8�~����~���Ͻ�?�м�U�A��P^b������$s	�e���G���W�ƍj�S�Xc�I�RE�l����-Aյ�9vQ�X_
+q�xۋg����Ŕ 6f���5�5�J��+��ɘOo_��)�w�����0Z�|%%�������(--�PJ{�lۋ��!�1$g\�4�*�E1f���uO���Ҳ*T��(3*���+��y�6T)낡���hQ~2O��H�s�"���f5��ֹ%>ƙ��ۋ_�Y+����n���*�'<���5�2591(.�&X�����~�
����qD����FYi7�5���ʛ���j����|�<K���	��*�98Ԕ/U�iH�&�Zy4�L��V�(#*'�[��i&��Ab��E��ň�AQ'��VM����h0*L�\׽f*�?���N1��Мd_��D�~����R>��5�Z-����~"q�,�����*��G�Y��W	�=ј�r��o\]ĕ�����#%�ۧ�j����\������Nq�;�+�k�^;x!��<b� ���w��FD�w���j��!�SJ!�S��&���p�\r��b�0r�8��F���p �̿P�Œ�}]��'�L�;�O�O^: E��2���s*��s��)3����3�"��R���aa�o=��X2�� !#�X陚r;B�c��ӭUZg��/J���~�������ij6]ۂK!~Ef߽�M�	���iF����i=ʕ�ŕ����F�O�r�!<(����F���Sr��Oѽ�>�W��g�TO�����x5� "��`�(k�ܸkj\��{��o�(�$z��#�����"���	qEP��z���^%�cx�L!�c�siǘ�SǑ���Z3��Fÿ�c��C��߾ye����ڎ�^�>�<:�߆R��2��q��k8?>�wc������?c��<���H�qT�[`4[�c�7��kq:^��!j�ݥV{?���I�|�
�y�mE���H��6J���P_%��R�E��ӣ^�I��uI����iҲ)��7u4���J�E��9�X��Z�TsL�����E�N�@V%�I��}�d���^�Ӝ=��(.����Yh?O�=��d	�z�[��'�%�8�<���6Yzz�KKG�2�ej%����Ĳ�P���A�S'���ރ?{�Z}�/n݊�z��]��XU���l�§w����]|lC��q>ea���rO_T&/E�s�{���|nZm\!��1X|'�Do��BAԍ���K9]�ɚfĸf8	���(oG�xnM�C�dM>R|G��4?���Qu#&���o]�v�Pщc ��{{ڕ?��ev�I�$Q��k�'��`��W^;$���߾s��MW��c��i7���tʹ�J-5;�8�k��eD%�0A�8��R p����o��]��z���ӆ���W�ʭĘ[�K'�֮&1>�R��M�P��s�����Y�WOH9�sA7z*�7�7����S����,~A9t�Q"�̸A���UI��Jaڔ����٩^|�|/+����m�老C�4��k���"�K6�:��p�iW��\�N�0���C9��h4gR��aNTR�OVc𬴰H\z���Qlo�뉦0���p���X\|!��_}�Q1|S1�޴	�����ӧ��W�Пb��B���t�)����z��t�*��2٣9��8Y<h�=�[4ZSb���F���/����h`�ɋg�Dw��Dx�| ������и��ƊM2�0]���0=� ������_�}5E''��G��C$�������防×��rv�����CI���58�(�_��w��>�DG�&Եl��dE�;���c2�L4%�󚼤���^F8��)�z� ���&��"����B�]��7���C�B��T��E5{��
e�"U�_�|�I��k�Veб�V��:����]Ės��Do��f��dF�-�O�&�u����=���XQ�Z�6m���'0��⥐V�M��*&�8X�z-g!e1����eI�?�m�]��[׈N�2])}Zd��cJ�3,O���k59�3�&#����5����7���/���^aƎۿ���v�DZ�������a0e�ج{����^�6u�m͍�E�H$��Q�����tm�7���ވ1�@��fl�D,��w��J�+���l��z�2��wN������)�͕I��*�m����������X[�߭�"�=(1FCQԖ;��c���þs�U�C��P�����TJ����醵X۽M��4.'����R�4Xp�vZ��bkV0:epV���nB�)���8hgl^)���Pj���ޡ���,:���[E$/r��Y��>���������Z����YPJ������|��볜��o�$� ��{q��p[������ee9Y%��c�*��
K�%�󘲜��l�PԠ�ݥ%�፼��UWUʿ��*yA1�Wv�Fc�	Ix�p�����7��VL������(���>"����S�L\񅋹�tZ3|�[��Y/��˹�C�tG�vx�.�}������`�
&F.a2�G0kE��{]+�V���a�����lZL��3n�\8�r�ҙ�bJ��Ă��،o+S���ݿN5Y�"a�N:$�&2�7ٰ
���}cH�,�eL:���u"����զ@C�n�	fd�Ǫ�{�N��������^�V�����*�W���ɬ��Š��Mba\�R�3�N�����7 !��:�^R������bV��ad�^J�+�`m�m�P/W>��6x��Mh�ڦĔ�M�Us��>�]T�i�Y�`*����ѳo!���~�t�����C����*1.-ګ�9�yCb����c8�����ء�'���)�c8E�3LQ��h����<?���=�L3;y��V�0�!�vI�O���L\Fe��0蹂��^<�U�����qb"cŭ�Q4�	��i3�\�9��.^�=e9+Mh�9�"�!�U�j�����տ7����\��l�t��X8��0j͞�ՋY�+rU}�.k8e���f)/]4���E��O(��:�� 8;g(WC�_ж���c��C'�F*q(Z�cN�x,7U�=}�	��?`�]�ȟ]��YJ����\�!�+��=��4��X��w���R�%#܎Y%�T���EKQhCX���O��i��.��u�Y�x_ؽAV
����B\����C/��T� 4O���h�Ӝ�N{ m��0�E���.�J�ˌ�	�3��+qE9B�T68�㯝x_��}��-����Eh���G�Lɂ�^�<�BWU%j6�d�"�����i�����n�p�Gz�j��� ��w0��8ӥ�E��sm�m�bE�g�g���I_�KKB1UeNĶ���a�'�W�Њ�Ez��v��+n�U����ӽ�pWJuű�	iN1���1Nhf
!�E� <ӏ�ou,^��� !�i6�5o��H(?�v�B{�^:t5�(�*϶��|[�!y�#b��Sk[i��'�i��б�&ɏPtf3�9�&L���_��I�ŗ0�:c�Ç��jl����؈HD�bd�Yk�n���=�3�r����Şz�rGs��CҴ�8o��������-�MR���֊���d�bc���6�uXR�"���K2��'r��,b����]�ޟ�K%�Y8A��o�;��3�;)3�=���n߈Dx������`$�eh�؂�u7�F�P���T�;D���OC���K��˥�A]�͂��0���Ӳ�J$a�|�� O��f�U �6d
���2��ě������]�]���|�Y�׭�4��C�&�mz��rg�nu�C�c��vIg������qɂ�r���Ȓ�<�9��]�B��`�=��$�&)l��BQϝȸ�VU!�bN%u��*ڱ���^ZC�K�B׮}��pZިt�1�n��5ɰ(�b�7o�,���К?Y*�r�\Y!�&�����7%��X��C�*"�-���C��ݒCg��rǽ��$�2@�bQ6�t�XGt(�}����,��)�3ׯG�R��!TF��RY��i�k�����_gBk@ �Ƽ�@��z�ח�"�P��� �A0�A$G�g�ZC8;�Q�����d� ����a�e0,�(T��7P%f�d�:�d�1rJひy9�2>�OO�j�35I�g�߫VL���@q�ʹ~I�2�lf�~8��׹E���\JWcؖA���6�D���S�b�(	�@]�"j�N[��;�o�,<��1<wb��E��AS�z��:�^\؋S�2��b��h���	�̿|�&��Tc���A,=����<j��H�ܪV_D�����B������!E�>��-x��9��bI�r*\8(J�r��i��+�qbԏP2+zc4�P�c ���}�e2�u�RY�FI��Ա=�R��狪kJW�ҝ��'����cM�w�N'*�|E�׺n�,q:�"v
�ѡ��?��_�T>DDq�D�o�����G��D�	'1|i/����R�Uۘ{��K�����s���B2�ŗ����L��F�P��TΣ?��Иbʬ��Z��U|�y�i1��������q��f\�g� r�R<�Y����JN[�6wwng�Ą��6��O���0)E<*�n��j���ܜGu��S.�JY[g�#MF\
��S)Ԋ���\��J��E���F�m �O���&8�͢�~_ޏ�}V�T��̎���������������P�I����9��:��QD�c-��ڍW/��̌��X�L�V����9��^���������+-xl��D���lbQ�~eĀs>,9(2���wYQ���t��:[���98G��ޅ̒"P:�յ?�aC�#���
��/�)�}<~�$Ք|�=\TFC���PրoxZ���6�_R��"��������U0L��1DS*�*�u�ƜU�/ˬ�� E1e����<���mk��)e���ӂ�λ�51�t;��J�e��Q^�Mq#?��u{O��u�c� U�3rGYu�Dte�u0Y�72��k��g�6�-��$�D<P ���"cJ��`��'˟XֹX��l��
u|�7u��b<`K5��`�&q^&�w�����)	�Lfl˴`[��.�hΈp�
�h���e$��iv�a͔�e�:򕔽��Q��2��t!�b��,e(svA_�LR�$K+��4�b�����QKiC��4��D-���q,w�Vu�f{]����)�({�r��G�asNnOF����=c^|9�|���hɂ�=��dMI�bFYok������~{���옪6^���W8N�l-W>;�|+�K��2exH���C�,�Ȝ�!:��>�L�O�3�ɔN(g�F!+��2HEF\���=W��
�������sq��e-q�7�[�#��ҥV�n�u��h��ԗ9LdK����倧L��1��a����2�D�dRQ�Ux���t��b�m�W��fK�&��1�8��)�E��L��R���3B�E��{�v�b[y��*e�*���rh�c����×�������M�T��hi�(u�Eɮ`m ����OH+v�]��!��Sk:�W+�L�R�{bnN&�G  ��҂�]h/t�f7��U�Õ#�4�嬕���&p�o���+G�1�)~�=���ʱ~���j�fC,��ӯ�y���p19ϦO���B��AX�a�n�)+�
3FKQ/,=��Qq��j!�Eq��:�^T�%�G6��UE���u��s��z,�z�#�q�7[��ժl�ڀu���>>c,�C����P��7�m��h����Ƕ*#���"FUZ�r��vJ)�{���U�Ol��~�X�)��9g�G2���R=��(��zh<�����V�U���uk�N���X|����Z������-[$V��&[����#�+Gwc6����_ ������ �&���x+Z5�-Z�6��в�5��������Z���k�.Jӛ2a$��ݛ���=p�l5���Q��%��KP�&���~�f1�mW���rJG~e��a����yv{#�\-��b�k��g����=un��͛��ы���S����]Ꙕ?���+����]����8�*�*�p��eƬR�.�o4[��=��I�,�b�Ty�~�����ֶ
��3�/�Đ[:�
�ۦ�ei��C�DH�'g�X,���aͦ0�G��Z��5c"
�3�����	\cv���h���h(l�\q�E'��4��R��$:��+%reT��b�7[$�+�My��P]Qt���!_�k�����ա5�O�:�p�[�L�/!��FB@�<3�7I��:5��q<���@L���K)��I1Eo�  ��ҙ����V����Dc�g�W=�U1٬<�d������5�2�l_.����b�I���L֢a`T�q&��9�,$��Br.��d�h�ٞ1���J�psG�o�;�?�����$j:� �S/�hV�'gf�&+�c�,��ݨp*g�l���
I)�=t� �$�ZC��QȦJF7�z�VJ>EY�J�&�N{��u�64��m��14(shp�t�@ ��b���i�6�J'�U�	�T��H<������Ԭ�xl�RXJ�i	��:W?���粪s�&�^���\�S�	ß��n��/U���èm�H/1�9̬W�{H�l�\x C�R��Q�B(9�,:6���)E��B述��.��pK�Q�����XSf��_V�.���L0�+O�f�&�#��Y/ȝ-��$6��)e�D� �a��� Y��[ެ��\,��!���RDLd���x��blԤ������;�+�d;Z���O0�Ƌ�Zt��`>���N���+��{�w�U��*ڷ�,r��W��=�mV�� �.�J�Mf%�|�%���i�(X�u33��B1B4� �/�h�w���d��WYd���Bf��b���#{����DFrKβ�������I"K`�����\ȿ{�0o�6?If�t��z�g�S���JY\�����<�@���ʷr�"E�86�i��~Ά.�������Vt�chS�#��2帐l`��:+�Ӊ��q�I��`x�d�^�թ�,3���o�>aN�Ъ1E�p*�౦�u���hn^�$�q���x�~,���C���G���$HC3+��8w�/SXg���}1���66�*���8L�D�������7��6���5űYD�s�l�Q0����.'����b˼"Kj�a�K/��H��ł�CO�c�ֺ���H���z��ڗ����T���͢T��V���4�
����^�+l��0��"�0�8�79�(wYar�Z���A� W������_�,ZƐf.��c��7�U(�����3��CgD�)�I�z�V�����rnqxQ[����us<V�L�Z�v2M��2«���˩q�qD����$����^��a��t$��LY�W1���a��J�h4��#�)����<�i1�!�>ZE���Q��#=�!�:ϼ��~�J���&��X�IӮ�¡�Щ%�� lo���8�tH9>�c���R�C߆�FҀ�L�pp�_���:��<
gU�����>�9�*����`C1�S��n���g[�|�-�}�e�q�b��o�?5�g��M���[1|r[w��|.�1f'�MY-O䃛S-Ҽ�Ǉu��y�b�G����H��^<X9��5%�q�?AYy�Е��c�]H��\L�q*^>U(Ǳ��GS�:�7�G8,F%YL�ߎw`�ĳx9\�Hƨ����۔�4]��KoD$kn>Ih����[�(�0K	e�_���]j-u:މ�/;���ŭ�V��H�=��b��$Ƶ.��a�=��5�	3_H�n���ـ���1yH�QR�2�P�- ���L�(����i�W��i3�A�P"��@���!�o^\���<�Z]����%���XY��"�2����R[�%�+`�N����1I�V�)��!�҈7ϭ�~p�@1UX�rg�������)�e�]���d�3�5(��8���L�_&VڌT߳���-ܚ�Rf<�(��Z5�E[$XW���h#	����b���4�Mݹq� α��Wvo���������J�Vo�}�a��"����:)�(��+� Բ��<��XDb�RR�غ?����y��������E�X�1��(�yA����`DĐ3�����D=�Fu���rH�ɮ�)�cO{�0����J#����C����+�,W���4T��Y�a��a�a"m�h�I�7i�����MI������S�K��Bk�#����c/�{�G�|Ӏ�ә4z/���Cx=R�X� ����n!pu�]�����3��J�'6
1)�v�℀{Ԭdn��'/���LtwL�*\m���{g�b�0Q,�  N\��7#5�P���йn�˵�	�w.�}�G��n�m.��D�*�n�A-���՝�v�F16ч��������F��P�ݻ'����ː�,���g��	e�P�g��Ր���@�.�UIk�+���UD��9���x�j[o�}��,�m�,�-]MJ�W�J9���>v�m'.)�A=�G�7�~��U4'���8w��;pCď��c�26�5�Bܮ�. �
 ����h�RC���aT߮�j'/EлWF�|�_�-�.�99�(��Wߠ��.1�	~��Z�:��URB�3@��	I���Jq �!���Bk@�g�Z�p�Y�b/̴�)��_��z�J���	��Ё+���͝~�]��J��±�N![��������CP-��s�]/ K��5��e@k̎YM/ւ�W���?�KϜb�}xLT����|�g�nEC���+���#�D�u��N]�Y�1�k��J|Ɠ�$p=��ްH��ݎ��_� q��4���kd�ټ[��߸��
x�bA��1��*�⌭+��! ����g�/�ļ���Bt���dawV2J���+�|����֞��r�U��Gʡ2,�8���#���Z�
�&���tKH�
!O���G�|׋�Nl��}x�ET<�͖�ͥ�X�"�t����f��觑Җ�6� ��պ�!ZY{eǴE�+�~�su�EY���Ν�������_2�q�0��ы�������-�8�S6�Vc e�_��78��u^{S;j�7H���3�}'�/�ꊡb]!2/N���\���>L8U�?y�]T)�7n�"���hFGk���xꩧ099Y�+++�����+�����׊"
���)��a��vE�ֹ�u]Ҳ���]����V��1��Q>���u��X��n��O���k�[7����0��㭈[������Q�a
���~�$�[)�a@�+�a�QS�S�\�R%3Μ9�o|��j������OJ�;�(����$�3�?�Ww��~z����Q�ǽ����(��i�i۶�]ߍ��a,m�p�D۾�'$Oo*������w�\��_������k8s"���O\�������7!7�J������7��p�����<��s���i��� )�ߵkWaW�k_'�A�yOO��_L�Bi��݂��� ⿵�4(f0��O�oS�6�_�^|?դ��z��:���V�ph���^��Z�R�o�iJc"o�^p��޶F`5�E���W�����آ�����?ceLd���������Y�W�փ|���H��z��>�\p�3���P�V#�8:�2�5JK�P�&{����@������g�ޥ�_��}�ӛ6J(��U����B�����Z���L�0�k_�ȼ�T(
_����c����
�4��b��@���MwJ��<+���Z�;4�.��_Af�-2�,�8g�`��}��0k�)�x��#<��GrR��DN�ʏ̤�cu-4�VV�Gd�eMUUUappp�UB��쿦��X��i	V+r����2�|!B��`E m���E�7��ꢕ��{�Tߍ��3�58��ح��{� ���V&������� .���G�l�b4dQ�,+�I؋���s�ќIg�}���Ʊ�v]�O_酻�_����eE�=���۽�J����!8iA����k���'j\k�Q�W����GM"-�˕�w�(��`��x�b���D)��a:�"�1%���hҢ��}��o2�����ۜ�̈́��v��!�1���AF�� |3{���K��|�wbxx?��ϋ�.z�M7݄G}t��^N��9/4a�i��J
���p���#��?���������(�ńcn��&�K�j	�=��+�D��S����T�n:��00&�d���XNށ&_uY��{�l�J��:�b=.��t���/~�6m¾}��U"&-+2Dg�jM�CYc@ 6=���6�/�Î�1���NEc)�r!jq�}�9��T��	wv���c�Z�g��2��fހ�5˝���lڞ�(fL�p�5߬��v�ک^����:Oz3�b��ly*�j���_���w%s��Ї���T��ճ������W@�7/��&q,}p1��\��p)O�"9C!�ϝi��hRΧ�݆b��Fl���G�-1#CY�|�����z�,c-d
V �����癎�.�j�Р3y`؋�}12\�GD��eq�(������~FciX�ׯ�[�����e�{���k�����<tn,��Pl~+IK�-�?�	����!��q���s��;s�Ϯ�Ϧ�!#�j-o/��h������X�$�x2��ϫ�N �\5�+�\�AQUmNcsIPk�)T�m.>�d�r�5�Ϲ��SiFUm�R�lLE��?��p��x0E	K,T�vK�e��P{��J�-&]w;Bx�r�5�p��H.�31��W���fAǘ������Ύ6l�� 셃�Y�x~�^EDY��lP'|hK���D��%��� �~�X�J�V�K�����c�l�|�7��E��>�����˰�8���lW֬IC����𣧺�ozTy�%���j{i�wo��X ��¥d�tԲ-����=tN���{�2�����۰I9�1	�j�KE��	���`ݖ{V��:l7_��~���1�v�:�rYc��e7JJ�H9ȁ����X�ؾm���'o���3e�"�VX���2a\����l�d���g��h���bM��m+��W���_�]U�ƶ-X��^�D��J��,�2�@��k{E&ZJ���FV汶�ag��������s$�m�H���9����r��S�3����)��S�^��}#J�����'t��� e~v[w��t3�����v�~q��m,�a�u���*�&7����G��a�6v�s�A�dLJ�gfO$��5r�#�Q[�1|��Q�ǐ��H4���p.n��.L�hF�6��k9��_�A��q�V��z�uf�'}��l��,Cs�!Tׯ��U��J���*Fч��	����K�İ*q ��г��܉��v�	E�>]|gGF�R�]�����u�q3�DH�_V��?<�ӣ��5���%m��^բ�����Ѳ�6T�DT�Cj���w��ρ�`������n��n�C1ČH<�s3~�kQ'���k���~ǉF{QE<s��:�1:JC�!�L[���6<��/�C8J�Z�0ǁH9�6	��HH�1�I�K�nͨd��()�<�
�K�5�����w������qZ��}2|//Eױ�_���ɒ�j�'#�:�,k�tw�bk�׫~ȼ��Ϩ�#�4B����y�P���K�tȒ�T	�S�n���Z�����c0��x�+�� =ߴ�:/CX}�'=��f�6������Q$n{y�ReW��d%C�+ѧ	c\j����]u�#�Cs
�?0�̸p��/��I�������)�Stڱ^�ڔ���Ѵ��iTd�Dz�w�It�J��,
E=8����I����x��P{$v��!�tf�^�g7���+�<u]��Gz���Ԇ�T������\.IIO�<x7h��z���aei�<s�Z�m�4�j;��F�h>�*j��⫞6x���£g����p�Qb4����uU�����d��L�E�:e��+�V���5�4~���[[�v�G�#C���Qye�\
���q�#�]l��pU��(9U�l��[>�\�	ܗ��?��e&0��ZV��3�ɖ�g�]T��2b�>�#S�zl�z��9X����8<8����詯V4|&���Q�nQ��$���)e���f�Eo)	�	���`V�s�ҎQɶu��g��4e�K�J�s;zP[Q��>���s��>c,�}\'����-є��V�c]]�c]I��w�b+���)"9�����B[�Nly�bHs�ؚXN��h1�����z��3�\n3�a� h,�
�MH���lҷ]�}p��}\�Pu�H����^p_���~TZ�(US�^���ze.�mya/��Ӝ �b��&nB)�Xt��F��2��c���}tk7+�d;;f����K��*!3�+fX&3���L���oՕ��ѮV����DJh�G4�GM�\ e�3V�
P�t��d9v�U��F��e��Ҕ3kfY�>|�(&ٳ��$jc�����L@�j��j���Ud
u(q$�5�
��9�8�؈C��5���^6qX�6�#A��W�/L��?ލ���ׇ�C?F���PQY�A�&b�=���O�P�@g�&��u��A�`�c����^���Ub
�zϟ�"M��[&�1\|�4^�Ԡsb �������y�^\9�*�Nx��g����X��e~=�F8�*]��(Mb����uXj�f'�^���;���6M�:�άNrj3�W�}�S$c��{G��g�zE�8�%�S8w�I_#>�;���O��Z�!��8.3���Eh?/��Hʆ��l��H��k9�9��DʬĒfMh���ݝ��
|�f\�k�St e p�]�RH�P�B6�B����ԗ���x��uY�F��+�`�W�\$�Ơ/�~oH۳o���"3������c���r���n��}U6���T���Pq�u���63�1�)�YՀ$��r�/R��n����F���
b
��}����3E�w����=���=������Ug��f�>V�)z;�}�]�����	q�Ãz[F�;����AUU��`�WOS^��~1C��ߢ���˽�a��mӰcF����������W��']>tt�@]�1{��!��ߋ�	F%����2�D�Q4&,���}����9�~�Lѻ 8	�=��s��{{���p/ܵ�b1z�.c�w�����jf��\NkKb��Ӌ�7<������ΟT�v��qo|C)��"������	�	7�g-����1�f�C�2�"�0��F�6u���Wr��Q�}����U� v��%�����^"\WV�"����$.U޺cf[�n��Mݲ�[$F�P���I��]��.�O�]%����G�/���V�b-ҊbY4f�c�L�m��Ռ���H��ַc�소���5w*4�r*��c��]Uׁ�5۰�wR�Q���Z�pմ���� =��
���*�	�%&T(���dW�)z�_{�����}��)�'|2I��[G�[w�D(�h�EHj5P�:����*��jE���\ e�����f: �t����V�d��W�u�&��ʠ���k�kYJ���},�)��?:~Q�x�R��p�O�Q�J�^H�-
ӛ����Ci;<��о�X,VI�phP���D"_����Vua2���X';~)��3���P�<��K� Lgr��r^�o��
oڌ����o�)�Ks������3R�5H�ݨ�'�Q~�5to�55�i�-�}g0pi�lJ�D�ָC��mM�:ᙖ�I��1CK0��A|า:��GtZZ���Xچ��8ۀ��(uh{{��I\<���{�?�2H�\z�߀ϞQ�\u�h�����˾R�:5hu1��YlM	G�Ɋ�E�Kuf0ӧ?Ňi,��,"S0�H�J��U�d_ĉ:s
�S/"0q	�V�;a�wx|O������^~p0Z!%�7G�hzC+&�b�z�"u�,b�u��Ŋ���|����)�=��� WY}M=��}QN+1Nѭ���l�N���A�@��|T�DZ10�3B'��Ja<k���-�Jʋ-+;h4i9�w���ae�>���y4z��s�11���t�A���e�(����U�<������Y}y��Kv����`�C��FUV��"ӽ}E�}B��E�ď�fdS�w�s3�j攼�c���!leЙ���7�!��U�f)��a�^h=��lX҆Zx(&d�7���|(��3c�b��+�G� P=�ݸ���  n(�������;�[��MӢ�������Tb�r��ʔ����J���0J�9!���!�'c]Zc�=�ϻ��U[����ط"�Ğ��x���K�ja���#���mqUH�;�}ؘ�Bf��/�z��dZ�~��\�נ��S����=��z�׀����l��W3�m؉��?���Bo�:����2Y��Oy�̷��mkĢ f"+�2`�ޒ����)+eFn����D���{�Cx��Ö���kg��l�����x�e��x����h�ޣ�Tg}�0�"(Ґؒ�Ծ��8n��	e���oym�l�@~����bʏ>xLY!3���o�*@��xR@A�����	���s�b�.�b�"d-J��ݬ$� n
��3��۔Ψi��٦�s�hn`U۴���i&��O=��-u�R�I�Bk���W����R>@L)2�^Ō���3�K[�X���D�͊ku�j�z���[��^Bܖ��ʎ��.�RLE�eD�ԇ5ϓ��+�u�w�m�h/�_V1�����1�*���a�\H&���{�}�M�s���܃�z��J��^�@;7W�FÅ���
x���$3�
@ʝM��7��wL���P���D{g�
S��L�r��KW;�����n� �$�g�
j�Mu|a�2ū��-s��+l����'�ҾY��ӆ>߄ )��g5 e�o�Z�"�X[�����T�o��f至��̠� �:�J�d�Ʉ-W�UӅچvT:5h�|΀��s�?����⹊�����j��c?C$8! �&�YjPG.��#�a�nՊ��=}E�M�sc>�2�=�	�_Ly����s���E�|����qSG��rz�'�B�u��߇�c��ҹ2�>�\9��}v�N�ϭ����@�rT��5�����$�S/Ë�VD������.��o�=�]o�\f胢�m	��5ؼd5͌�����&�5�&*�F�N'���Q7�F\�#9�J�Ͱ��N٬�����������h�J��bJ^K\_f��Qס�F��Y4g���xY�n����Wy�y
g�N��^\  ���Xm����y혱����9�T,��~E@��;H�j1�:3c���� �l^�y�㑿>u��k͔9̸~(z}�NI��`) e������4�Ld삊Q
}��Ҷ�˯.Nֵb���2�̔�[u�x!��@�z͆,�Q��]�?����4�\u�[t(�Ao`�q.>��A�V�����c��^�r��KpS���|c� 3z�Q<\9�.W)\�	�x��8����&�xF�!�d�<��oh�Ɔ]�D��^�v��ϼ��3���Vi�b�Hn�F��C�־�Ɠ<�\'fX��y��fIK\�q|x�m�%��Al\�k�܋{��;����Qz�"��i+��Y,���̇�UVl��s��V�5��;>�t2�{��V��ɔPC'��!+��w�I�*x��u�������$�:���R��n Ʋ����a�[>���l�����'���R���F4�-���z�zz[4�c��u;en�Bْ��E���5h�]����1����+����7K���d�O�� �!S�
+e1�\g�a�}Qr�X��ڥT WHc�N-��� Rv���ܱ�_�[�*�ܬ�|�p�j9U����p��  ���[L��R9>4�-M��%����u��]�)י���\���A�I�@k�)��IH;�z:�k�^�0�(��A�E0�Pp�h�d��Q����2��M��>�c��pT�Ο��#� �|\7p̅��~XSm�_4!�V^���!�0!��#�@MC�\�(�#�5
�r��k�L�R�5&'v��T_�o�a�D"���p)nC Ch�,܎������H���1�ܯ���=5[��i+@ʷL)S����4m	�\ӸN�[S�Q���p�1�G�<(�@S�`̉��l�A��{�j*����/��P��l��|Ѹ��L��2|F;��^�)j�����-�]w?������!��kCO��|(Ë�Zt��`�����,?%���g_�O�b�s��Y����Y9���~�r����h �C<�Wr���j�ӓ�K��c ��x߰|ɔ�ĝ�ȗ;�;�"i�-�C�ۗ����4$�Pʆoy[�k��]8�"�B���mx6�,�7���$�e��e���≩�0�q�7�@,k@sIF�����D?��쉬p�o��7:#��a�ro��h�ڬZ�e)}1�n�BkmK�����<��^:�l`U�'�e0?@"����4�>�yL�D9�L�^�D�5�?Ĝ_Ӿ�_�1U���h/����A_�Zl�'g�Oۛ���lnVG3�]=�i5FV�$��U������w�h�9����^=|C�q�)+���ņ�-�,�d
��\ح��.�zx��\�T~v�Y�1@���Jv�R~�Ý{�񦲹U	����aS��ɀ�Ю���_�Y��ϸ��2Y����������4|B��.SJ�Ɍ���5o�PJ���
�8|������R<+��@�,��̠i�Ж5bY�y��Y���c
I#����o�gv�`\9��D��"h6��c�ϟ�'G<�_r���7H�ڲR<����?E�]e)��=�����¿��ݲ��~�Ox����n�G���l>K��cI���	�yT��Ns�W�csi.G�L�qe8�v�Hu�wCx�5�{�S��t�rd���!�:i?����uO�Xb���o���������.�޽Hp1���R�Yf�"K-f1_8{��_�=i8p�r�t�a�����A�L��g�T^r3���}�������g�c��~z�����=x����qebS�2y���t	���s;�_��Ƕ7�n}��&���;��c/�=4"!x]�C�Й۝1l��WP���e(B��^��JW^��MN���F9�;�<�k��.�8tfI�K����V����}xt�Z����⿾�_v��$�'���Aʵ��:��C��b��f�6�Lf�y�"�y�W��uRA��}�y�w�n� ��}�L.yø�9�͵e�q�a�W�5�7����W��A�WNE{9	����Բ5��;J*e!��	�۱�vl�>^g5�ey3LPj��1����YN4��M]�Pb�[����[wsG�݊\!,I��O���Z�+�O�{{�%w�
C��t4�5�O��m�2�o��"���:��^EO�N\���cS�;�3���XB뚏�TMl��+a(��:�5��މ���q<�!����-�p5ʇ����YlMX�,W��e?�@�(������K�{��7�yÄ�����E\ڄ('����ch@Z���b3��x!mWh�� �x<���ާ��-������T�g�WW�Gz�0����_Zp�P1�	J1L����58uɇr%��uT$]u�0V��a���ڒ'R�T*,�I�Y�=���˙�LƑfy��2)nnh����]yp��y��V��iI�۲%���q0`;�i!G���t�L��@�N;�%%L�@��@���f:@&!)�6q�����6�2�й��]+�n����Z����dO�̼��c�����}��}^�H�t��}�,Pm$o~E��%�����*���7�:��^������"H}�]�{��Ú-�<�3�㟞8�}�5���3"��x}��.���n!ru�-��?�S��M�zev�M/�a��k�%j�]8ٺї����Z�i��NV*���Bw�����,�~�v�,�O�[�C����rh�a�������B�V���(�-�<f�&���/�w1BbS[U���a%n}g�(@��e���4ʗ�ӠE ���\��|���B���^v�6"���Q�����+�}>\�{M'ph��~��+�\*��y���[�������b�EJ1�:����,�,ǉ+�
���^β3�Ch��&��ơʾ��*@�r�#r��>8�k�Z�99y�ۑ�a4|�&���B��3C�N�b�9�bܭ8Ϡ[4�j�:�v��݆���p�_�5ř�rn*����ht��f�+6W�bIp]�>�,������g�:<&06A� �ٽ�v�#J�����ӱ���wM�8�Q�U"��xZ��y7�=�l��5܅~{&��\�\�W���#8�Q���B5zcg�ZW�s�z�_��{:���:ԋ6�����;��{���7���w �r�+X��/�`�E�PN0�߆Q�Y��WcLQ�^��Jۧ�Vb�� Vt�W#�s"'G��8�����]����F�����VWh}��m���aDb$#H h\$���AW���i�Є=jq���)�z9zO&k}F��L��v��|ۤ�Π�#�$8ۤ��	vr3�6�)8+g���L�Sv�o�r�U�2��͡B\�R��u�[��}981�R�턅�iο1\,+oeD�"�D��j"<��ن�r�<9.Z�U�HR󍩬�T�9�G8q4��f�>4�S$��b�G�wR���:�o�9��n���q�L4�����H搴�F���H��#GT7�}V �@���k�d
�����Ao�\zT��TK��u�E������T���M��x�����M�[�'UO���Z)��#�S���s~�(�4�>�ͮ�l\6��.�i8�ܨF�9&��=��Ry!5Ւ�Z�=%=^� �)����י�"\���o���<:Yg�>�s���W{���*�2��8�Ӫ2�h?���oFIf���Z��}���`��E��qP5���A,Ms@�a��{0*�(O����E_?nط;�l���-�e��&����kIi�=���"�o�B�G���xщCf�r@���R�0��FM����AeƘ�8��;>����p��k�sE.�D'#
;�{/�\�I�f�%�ıX`wd਌�sԡ&d?�Q(Hs�\��ъlȹ2�jeВ6~��=K�C�}�Eؾs'��b+���L�R���̬l�9�Q,�� ��L�/*4��
��.�2kw� vd��(ï���q�x���x�ָ*w �����kP�|c��F3�\<�U�#�i��\�1nپ6윫))��E�Ox�v���!-��x�	��L�b�֭ؾ}���s ����&��1�q��������yΌ�ЫLی��P5��B7��F��f�ʬ!��Ƕ��nkYی���Q|��[�]����Z�Ҫ�B�M�~�>1�����|����-M������S�`�`�ħ��f�o�EŒ���]�|2z����>��]}ʖֆ���t5o���՚}Y�Kk|����k�j1�G�N0�WqVo��_�1o!|"4��Ng
Y�I�/�.����l$�b4��EK�'�#��k�u�:s��.mt.�Z[S�]�b�,�^Zc�cT��n�YZ�k�]��D��u��/�J]��)��ʠL]'�6'g���f�/-<#��k�n�P��-h��ҌI�2����1� 7�5���ԍ�Y��yvfi5C	 3�6��KFF7��[V�d�²g��Tx��E �eɣa��'1���/n��ӷ݈o���ۚ�:e�-�sm�ǓV�5���Bog�R&�2���NR��v7�w̯ˤ�b���sZ�@�9��U�A�� �%!�3�m���|��'�H�Bn�DB�Dӻ��5P�(3����6��5�*���׭�ҍ��p��24v��V/2c��Ԭ* ^�w�\�ϾHo/z��5:��_wT��n��WX���v�7���Q��z{�ƾg���1��=q�=��Cݓ�B��r��p%� CCC8r��H_h���뮻�m䄑d �� ��7(#���L��*���m�H�� 5B�$�
^��O�ѵ�WlVe����4�?�����IT���������w�Wym����'�۞4+AYn����~]���z����Z���mx������ۃ�JY!{r��46����e��|�ǲ����-����5!#X�k6W���{��U{Y�������D��!x�%t]D~Q��Ɓ���������ٱ��oʏ;'3p���M��K�;aӍs�����ܰ�
?<|R�X�0˩��(��%PQi4Ӊ�0QD�����0�XH0�y�����ڼFӔ ���s(�3j�KOl<׻����[W�Ye�n������fx{y���\݄�SqDL|_��o��sǽ�n�6��Ki�R����*锠�	뤪��>�X� ��6�+��fK�E 9.�z���;�ke�it[�_`��.Բ��i~=��HlRo���r��ru����=��[�7�0�m��|h8�`��H ������2��<I��^�����XV&�J �/�z�E��[�S؍g$a
3)a���H���'�/�s5��ʤ�� ^��!a�]���"��V��
T� �#�z���% ��Du��F�d�&qQW6�K�{�E�₨y:[��3�����B0�z�!�P��� �^FPÞq�k�c[�Pf�
)7�rpz�`Fɒi��j�n-lEma��V��æ�-]㥁2�X���R�}�zT��i���n8E5d�U���3����`6]c����|Q��������VC��G������.���d�>���gݍx��MbrLS{��}RKkl_�v܄�lk�h@L��~���j!3�"���t�_W����;���z����m��ΡT�N�[�@}bX����K�l��:�^��vj�O����!8N��tUn*�C�w`wv֔`��k�������r�U���3ޓ��h�Kg.���R����7C�k�a
It��縃A�	)�Iy�TS�d"Y3��ŀٟۅ+6�f�^���
!B�:��|=������W�{�9aK}�se�v�����`����%�NTTo���C�}=��A�DL����74-�0��Αe����֖�x�=SVV6g�6���������؍�(��`�s�U����>�A���YT,�6��_M�,MG��cˑ.1Y\�l�Ṕ[��O���ە =�Q��z��&պX�YB�ܱc����̍R����?����9�R��"��7��kBc�I�P��|��Չ̴����)�A-�^܁�63�W�HY�7�v2շheR&03�������q�2;�/�\��9s=�DH%�����i$>�cP 3eܖ�p;�V�V�L�-���nF�d�&�O���Jw=�ZΣ��YY��0��wF�����Hvh]\@�Y�s�F�.����R�Ő!LP�%qg��9m�����aY\7��e���E���安"�!ZVk��85Z���2���� ���E��d:���A�#8�хׇ��!хr�z�?�/�r���J�BP�D���k�T��L�����.J���qR���P	V:��v�'��݃��%mm�������[2��)�}�'{���:�d�م�fp���/��]��ﵩ������d�7j\�L� _�J
����Qcb��3�lj���9�<&ˊ�l��T�l2@A����̜��4Y�6`������I�YK�]Q���Ƣ<�ٿ�T��N��_�J��4���������a� t���/Kq�[�2.���;Y��#<���{�~�ӛ0>a�y��Td;�� +\DxAD�Ud���M�R0����ĉ*�w�ܩ�&2��=�v�
�6��� VMM���oM�y� >�����ǯ����:|���زe**� �566��߰aCX{��*ǁ}�9q�]�c���*��[dG$>~*�C��N8��e�S.�&�;�f�G򔘅�i��O:�ʋO�G����ÿ�g�j��OW���E��*�(
%�Ya���>��F�~�i��W��v���Q��3Ϡ��ZG/�O$S�]�jՌ٣�a�����E�����+���{�w�y�>����s����#�<&��3+K�9�
a�3ٰ�<|���^�||8�5�}?`Ǆ��,�>R/��5<������9b���3!(3ΰ�HDr�e��8Z��y��D��bB`Xg����oy-���<�\���^��Au���Α���$\�4����	`#�KKK��k��"	����=/��,�/.AX�Y]eX ��&��`TY�611!p�� $�\�9>9�;�Qc)�uC,D�F�w���E�ji_���ٳ��`�'#�˄	ΐO��g�<#�Ҙ�E�o����E�M��J�S`�8#�/�} �I\"0�^*�====J�� Fsf���ҫ�B���_2'#	B�ub�f&�Է<%�Fi7�G�2��U�q�'�v�?���%��A[HY��#J\��4f�S4L#�+�:ǐ�L�0������o�|�D�قU�`\g		���$��\	b�?��Y���c��O���Q>V�vg7e
q'�G�c��Ĉ��k��i���\\� Dp*�=409�LZ�%�f�7����ރ��@o4DD���y�������+i᧕�G�q�'�C�K΢&Z��O��!̖���AZ�-����px}�}#�]�h�z9�YI'��MZ*��\��1�O�����>ĭ�aB�FsI�U���7<����yi���j!M���u*��E6w���ۤ� �E�Q�e�|�9�V{�!����4Ї"��%p�����1���)0�4�=%��+H�Hgc<0�ԜU���(���Xn�q��v��r�$@�='���H~�+�lND"�'��#o�e~E�-���{�X���؈(q-cL�]��^��Ƅ|��n�M�6�3��X(��+���3����E?��W[[���v�]�vzDOڐШe<�Dc}���oN�(��c��N0� �`�s-,v5�Dx�v���<�܍�[Y�!�hd���y�*q�1G�ƍ��SO���qMΐhGd,0���&Hy?�����~;n������}��:��t�k�g�)-C��M��
��$+fG|~W�s�?�2�"](��D�K��"�"'A��TҀ�}�QC��^Þ={�nݺ0q�	�o)�r~$}��n���ٌ����a����@��ov>�i��'&�ym�jݸΖW_}5&["AȊ�ĸ�٢�]]]��r���+�����L�;v�y6+=��|����('7mX�����Hnmm����!rA�DC5�j,^knn��Ç5J/�n��__�L�M���xg@��|����/��X����=p� �x�pNs/y5��"�Sq��]���E ;�]�w�x��򗿜�pT#4=���g��-W��x����g?�H��U�b�_ ��y~~~~R�׬ĺ�k4Vnf �tP�Z�f��p�'J7����� ��rd߾}ػw�a$�wܡ�Rq����~���l�-�ܢ-:�$\���j�����&OG���O����p�f�\"���/3�J�Kau�e ����$�]�,�^���*�,2H��o]��.���)�xH�X>��]�f�*E�P16�X���C޿"    IEND�B`�PK   �D�X���(5  #5  /   images/50d22222-f918-4c14-b9d3-6f9cf2edfac2.png#5�ʉPNG

   IHDR   d   T   t���   	pHYs  N  N���   tEXtSoftware www.inkscape.org��<  4�IDATx��}�\ŕ�y��t�LO�9�F9KI����k��������~��p�w l��L!		�,M��S��t��ߪ�	�F`��ò.�t����ի[��snݪ����o��S$�R�kY��VA@��O
"V3 �����R8l�d@G���z����c*�vjzDѺ]��LA*C$���)�=}�O��Ĉ�C��4��=�zED�qz�1!��k/�4� {���4���͓�f�:�*�n����e�Wjpq|��m��U7؋����0��e��y=UŕhByQ:'F !G�3��q�.��ݍΧG������׮�	����FD~�R,�\���� +�02�|B�YʺpA����D[�>�bG�2ȩ~}l��T�8%k�KQD�
�B8�ێ��P�_~���ʦa���C7	KK��ݟ���7\���>��j���[�ǉ��x�\`H���6l�X�!��T.W�?n�~RZ\<��P�������������9�I���x[��<~�BhP��o�LE�!)!�!��|�y���_� uXnb2R)&�||��W���D����\�W��Dh�KE<q���k2�������w���-;ހ���IR
j2�pϲ�$�Ǚz�c���9��݂��؀�]��{����m�����I���w�mlZ�����߻��*+Dm-��T���_\�cbm~	Z��7���m��w�R��ol��5����Bɏ��@�ҳ�5���O��N�r9��/a��$m&�\5��6� u���4�`-j�읠�+az���%��ΕI$x��q<t�}x��~J�|������U�;��������/Tyo�����B�Z&G����	-�E���}�D�Ý���'bEN7)��Lr��v>��#8��I��:�hƛ�O#�n��=�z֩�8�&�_l���K�ɿ��$�Mt���2�/ԝF)��4�0/���kOBI����oc}A�$��O�ف.��do�55��Gp��2J��h�{���������FAR*��s�ة�8#tQg�1A��}ku~'���x��Y�-����r��~�����a��  ��
CO��/��bb���{�is�tM����4������.��UT�[$pv����.������%Z�0[ޛ@�aGh�}�ƻ� gz�li�Z�W>�5�ɱ���O`a��6�]G�w�q�����w�tO��=gn=���[暞��	}�{.`yo�j"�YH����<��.��*R���+��/���]	�B^^��ű�V$���dj($rx���C�(����n�R ��zr�I��̠��������)��D���4b�����K��7!����P�G��k<D�Bd�$�+�߼�y�b��%�JR��4�D̟X �$<�cG�do��[yoE�{�J�u�����8�كSx�#�3�]��A_ ֈ}w�P�q,t�cՐ����H@�&�n�"�*�Hd֠L3w~L���͇�Ͼ~����2���0�zc��Ÿ}t&�&!'#�a~�H!C���@EC2鄍��u��~�Pj��ϴURBb�42�~NaǤrb��D��V3�ˢ�	��~㵧�4:�����+��Ӊ��c��=�������BiIo�Ų�t,^����1,�*B������=r��������+������� �\�GO �#��َ�����q��ȴ_�p=~{� �6\N,%,L������wFҖ�8�-���8�sn�:���%x�;$ABmb+:�,4���Z�D���	-"⏠@xV��#-ƥ��4 N�?�	�!i��\�x��_�MlD�Glf���K���$�ݼ��_ +!	�|'��H��u���& 	FU.D���2��4W�LY�"����&�Z��c����_{�Y$�����a��1�0A%"�����HK;�_�s�q����IC9��GD�{o��/�j���u��eH�.��GWW���3�`�C�{9��QW[���<x���)�����آV���"��+Sq1ߎs��w	$��4��?�o *�9�T��i�\G	r�%�� �8?_N ��N�mr��ok���#���׷܌�=�ĺ㰱j%?��@n]��[w`hh^�7��	&w�Ņ��r�{�e�V���D���?B�gV縰u�b�F�+1����8Wv��ZHER����%���u&%�!B�64��<��IJ��fE�Dt�eBI���CN%��x,��p�Gow�����wO� ����"�8���)h� �6�<h��0��rHZ4��῵�3�����ҡ�*1��`)B�Z!��0G��� 7[�@t
c���IH�%`�ʆ�ϾE�ٌ������۠�񦞊�'��c�M��z#\����K��Z6E�<0��h]��Z	)���(p3>���Ġ�㶚��{01e�7�\F�RƭU�!�1���~DD��m>.�<��AP�'G��=E�$Byz&L#��k���9)��KF8(��'��S偠�yf�O�(
�������n�p� ���̏�X�L,��烄���&\[��R���,OE��5�fN��
T(���@S�o/	��P�a2�q��1�ر;/�BX�V�WT&	{��(UXUXΧC�Sg-���%�E"AD؄>_����j��_�~|T�@�"�gNU*��!a�ʔ4@���d���k����'���F�A�P�% �Q~��=1	6�n�#=U�`P�#B��iÏ��,T29�I���}�cu�
�a�h
b��P��=�xH�#���O��t �� a�[����"	� �	�B�<��"�b����%� VF).��R��.Dww/g�yy9�k��g�A9�gFȋP=�^�aQ�'�L�Dd�'"H'����Q�2�
� �sB]����NMa��U���z��L,��X���U>���b�>����|�#&qwr����d)�8�zQ&_��;�� I��̺4>>�ґdh�*N,� �2=p,��tw>�q$���JhU:��}�~͡�6�J`�`o[ʈ ���4<�{����(�2x�ϟEzz�%B�0Gɻ�R!Ab��F7���ذ4��`��.b��CC��s�k˂q�~�
� �׃T��	w�u� �H 0J c�;������G�6�E����~� ��OR_JQ�t�)0Z|0��m$�}�,BYr9�n'����xa�n(�AHe"LLNr�D�,�J�ӑGC}?=�=<M'ޭ��I5�c�����������V^C]D��	˴+��ķ����LP̈́Q�7?z ��Bcr�2��_��;Ӣ!<��Db	�
p
C�SBu$_J"$r�U�9H����@7�w2�d�h�Z�	+�"£� ..	i*tvt�NW�p����}���H�Q��G�Ƣ�*�}6����9� �K���|�I�=���pX�_��ZOs"�K���T�?�=
)��p�1�҅��k�+`�2����yĒ�����w6)ihTJ��jtt�0�f�jw䘺*ۋ�P_�̤�:���/
AۖH�_=�z�%2G��?��:<�O>�X�Z|�|q~<��X�d#&'�1er�pq�e_t��N����-R��E��1x�\e�� #�Â�:4Z�y��=��|hj9���. ?�	�JǊ�s��qEW2OC��jS�E�q�6",��5����9�[Kqx��A�J�n:��eg�DE�"9� ����e�x�IXִA<��GC$(�ƏsYT|��M>�|)l�A���ԽQ��	�e����7M�\"}�ŏ,A�\
u��ˋ���Ln>���v�V�%��p���}�.�����-�DH��O��g�̄�syQ�G�T6I-�{X��A��� �U�;�.�(�"e���j>u+&������Bai���K�o(i�y=HUdއ���b~u�M"��)#j>V������xT+j�=��%�>e�r��v�i:�a� ֬ـʺ�����K�J�X&����\qŞF/ҺVa�:���ݟ���06:�YZ^����z�;{�[�)�4:qC�	�}��M�D��!�Dad��t���Ƙ�+t�FB�r�E�R�/R�h��4��6�R�I��My�(L�J$�%��(/3am$��ٲ	]�p�ۦ'�	,''$�[7݊O?�3��J�?�S�v��Hy����&l���W���O��p���R"W��Fb|e���e� �9�s��5�1	A"�<G�^.e�E���?���]&
����0ϊ�%���;�4*V�od�L�r�8&��o�o�86��k7ޅ�����8=�K�������dv�y�л��L��R������㥪y"4�,3HCJZ�1����k�t��p{�R��SA���,�)R"�n���Y3Y�N��t��"'�Z�2`2�Š�1SG�D�r��^���S�����Ku�B,��:�<qFl^�~N��&�#���
��]����<���d�|���SX�$H�">>		���i��{K�KB'�t���� ��j�YL�ʱ���E ]=�g�(��
m
nH���G���0��b)nM.�N"���a�y��J5H+C�Ǌ_������$�RJ��gڻ9!�����4��i��dB�J)����p�2@�����r�wL�������qɸ7�����o|6�e�陝Y��"∩���\�(I~ ߪ+J����Ѻ��ʑ��Vj8yބ��������aWoUE�YD~7 őu0Y�taKY��a&�pWO�$)&"�0����QY �ː����T���p��5�ü~�I�1���d;��l߱A�St�>5���(�_m�q��{%	m�do�ۋ��
,]����T�R�_�@sm-6n��ڏ>�6հ9�)�M7��	o�M��^x}?�[���#�H��7��sx���rE>=�0����7.E(7�;q;Ї������o+�sҌde�U9��#���H��3����y+�Bu,�O@Yן�}StQ�C��k��P�� �Q␤>^��H�ح���zit��.<q�M�.�(J�,����A�r�D5��s�p����D6�.ơ�~�4�����k�$D�����#��R�RX�����]���$!A�$_�(^~qF[#dw3�q8߀�����RR��"9��gc*��N#�/�y���]��Mu8���o���]�%Ӓ��bx��j�B�qU�HTǡypͣ��O���a>�k�sK'�x�9��Q��c�(�-y��J��#n_%u�0?��ݶx5�7!L�6v�:�brf,�W?����.j�8����9I�qHJK�B��I�bB�<���_�:�=��|�J�Q�C�ݮ�ϮOa��*��.Ɯ�(�r,��4@���z*亍<l��S)X�4��2q��:���"��ƙ�F��(H�pv�#��L"�6^�S}AGFy�/�L�F�Ƒ�]�2g��"DӘ���s�v�%�q������녇x�Yj�::���~��Z*B(��N*��9v������.vb��s�%~��{�;\�i�=>j�4:�����	�^ B�N�����e�.4=k[v�`������F��N���~���+�;��g�'�xHfn�ϜGK�$��	����ed�S�Ƈ�Lk��|��皮�&O�P�p�>�%��?�P��,(�+�R���%pdڮ�\�M��6 �^_�r3�M��Eh��U\�j35Ϟ9�m��/F�e$�9d%='��k�òd�s�b;F��g��f���S?��H���a�6��p8�y�;7[��N�F��l1[B]7ԋ����Jl.�BEZ�4qh!���f���^s-_U|�9���c�:3�7�(�&�ߜ< ��������O��z�>�´`���p:�� �����ｽ�D�PSS���:.vs����j444�������y��f�J�D��a�s�Ш��^r�v'Y����RI�9<��Ij�7�-�S�ⶪ�8��A|$5mB,3��U�c��^���d>y�Io.�����rBI��K7��G�qb�����|l��v|b�o��}���#��z�/��2��N. 6���ݍ�۷s�G��i��d#G�3g��L�!~2�LPW$����t/r�� ��#Α��#A�F$Q�P�gT��C#Kg��܊)������)D����;!$�% ��K)��4
�-4�5*j�V$�:����㱚�ڃ{��Óg��n��q:|c/�i�eg "�w��X��$R"	�>��u��f���F?����~n���������@.�#99���� �����i����w�/�g�Mwh}�~�iI�8�<�� j�.���A�RȐv��(,A�(�3U�u�Bp��<ݯT���B�;�_m��5z�M@�T�G$�A\�mDez6��XGN*')���XVN��ɉ��L�w��̒�����iɾ}����ȵ�b�pM`����099�}�&�i����:�e~DI��1�b�Nrn�2�p�U�T	S��y2��	&�:� ���
�E��@{4��u���j�WF֦15��C'�T��@��.",���H �f�_|�	ށ���H��"��o��g5E����eAW��Px�!^�0mc�:]�:�������{9�����N1�����M�Ń��Ύ33u�di���+$ۯ�'�.���i�+�L,�����ɮ~���R*�_.��׫�/�ٍS��P[
F�}z�w:7�e�al|U����"<nÄ�H�$bBl7��9����± �52Y���t��ʲ�6��`ɺ5�ݮ�Ĳ��a�v�� �`��s����������1h�fv�^4Ov��������u��9�3�f�`fH+���v b��a�	&�A�Gf[�R'	��x��DX*i��o��֭���f�V��}���4#$#S�!3���001��[���s�	���..Y
�	�+9����P��|�!�Bݔ�4&^��5&�$�����F��P���	YD�(�/D~F&<d�;۹�_\Q�}+V��-�܄,-���!�r�<��mHKME��V�2�~q�CC(+)A�!������u�\XZU�De4�7�q���V�ZRV%�ZV���ڨ-YԮ�<HEb4vu`xl�B6:a�g�@D���$C�~6�t��pM�"�n�jLL&)]"F{G;N�>��/��b�1��j4fa�I5��� @�=�H�#�X�e'vV-�ˬ�/lÖ�}�{��ͩ����.�� --�����F`"9u)��8uz����t�$����_���!��pr.ҥC'��w#�0�E�3��W�����y���$�	!x7�K.�˦>썣{�%�Ylǧ�iX�M�/G[К&#���6��ӹ&��5 K��w�X،/�V��e��RB��Tw ~�w��
��@,F7�����P�E�N=��tP���"xKG'��
9�nO4B.�j�U����s+	�z'��]vؾR{Z��8��lی����{�kPa��)	ص�Ɨ��[��@��)XB>t��Ѱ������ �4�`s!���y�xq��O"�����ii"�-"!���HlE+�SG���q���G�i�,t��~^��>O�=��OT������a�:�_=��w��^�X����\*B�1|&f�Ȃ���+@V�ǡkh����aCz	���,b&�����H�㾋�:6233��pN>��[Ըɛ�Ǚ:SW*aҒ�J�j�XIN������ϸKw��C���?{�=4�{<�;	3�YGD?����<r�q��-C�d��޻H�]lV𒺁s��+��P�G��W�a����r
�>#!�d,�H����h �Vx,.�M| ?=���M��9�q����j)	QF�n
��!`�՚ ��O�$����(/-��B���<��!Ԅ��F�2͒`�Y��~Cd���^�+/���&7��!��Kj9��g�d���n�4�������w������)l-߆�q��!$˲�>���	�;i�nW���eS�8����x�W��Y�'K����6
{�	�<sޥ�B����۫��_q^��>��D'4�	�+I@;
�hdЃ���F�P��*4d!�)���;u��t��1�̨e~�����X��+�"K��a�˪��^v�[$y�X�?K0܇՛n���*�Zh�:�9����So#��Hߩ��8��'j�S����>W�����.,��N�lz{�w"��T����i�*��H,������\�&��5FH4�0�F	� q�����/.�'�{��]�y�N�h���蛚Ċ�B���P�����-נ��x�Bzmw���R���/R�+�ੳGhT$G#���G��z3�4�wt(�W�̴Y�t���e���ۯ���ߨ3U*5���<�vt�N��I`A�(��;�>wt/>��&LC��i���I�O�¶�Ex�MK3�5��3Sp�.v<�<�m������N�!Fn���>����3�.����29�������脣��Èx(E�V�d{F�:5|w��9�/���Vm�7w?�kK*��,���?dǨ�3+�KR�"X��G@��(�q�=��ض�+�ę�X���w�d[K0 �b�i|����W��b1�9wU�8�ہ��q<��_��T�	��D�X��w�#�۾��N��Ï>v?^i8��݊��6�����K�l�����g�[�G��>�Yi��1�a����+6�_�m5�x�����'�Z�P�R>���e؇q����g32^����6Z�sEf��0�C��!�;���5�;�����K�Db]6�|�ȴb�k	a9�>��c/�2_Dbs�)鼓���i^a)1�'N��4��^&�����2�N��踓CΈV�*D��ana11Y}?��>�r��;I�;����[K�d��@$�mRp�u�2�-XW��dO��.�7Cvlߐ �!|^��"ʞ�����K1�$�����m�<K�<-�V-e�����8���we�W*��}oĳ�O�7w��څ�n��[f�sח/���&�Mz�L6�1�kä�w�Ή [�D���*��Jݙ�*܀ ÿ����rH�}%�f��w���O����4��F�֞Cuu2�s�I�k��\�(��F��w8�����,Ŧ6�q*]<���.�e(c�x>�
�.���l� `Z�:a��d�f�|S��.��������n���NZ� ����5E|b�m�����˖i��ga{�n��=_{�/û@b� i4�g`�Dyd/Z	56�p��������}疏��F�\��Wn�f�7�]�
�|�l���͙]T���3�󄥜������ǆ�O���*\S
�����e���@��z����y����5۬8v�v��Ύ�����/��%A��4����v�n�?H�T�cjCgj��A�SF��'��eN]BN�?�)���"��N����[<p�"��=q?~�U:_��g�y3��6)��1�a����=A������e�"2�y��<�Sv��V�����^/ן�{�2a15D������v�l���⃀������`�{���af{��g�%����ᨯ��jIZ⡠ 5i����F��(�7o�pG5P �����U�����0��{ںs�&�X:=U�V�*Èа'[]F���^&Q�=�d2��e'�4:��ZGm;olei"������3�ԏ	\N��E�=u�h�A��v��Q�W�7�M7��=��V�}^�`�� 	t�j�AS�4���I�Lv[�9�fꞾ'�G��o�b��.)�0-h�x��,�'�CGlNHN��@�Y�'�*�4'|�bMM1��zx����`�7���O���(���$��n��2A�s���Bj2r�J�&R�[�����|3�;��Ɖ�14"sb���\��\X*�|���=~�G�,+�*�[�\;
O����/�%��AY��3�[� ��$�@�@1�
뤑3�g�0?�]������(�\��>�渢�pO�r��U���8TUU�yqx!�4l=ڷ�`��@Ύ��}�Y~�����N���%x����Dzy	�G�b|�E�pB��CyM5"���$�9I5=0�r�w���M[�s��GuNSo�#۰��0�`!ӥ�5I_��f5�w�#����F0�N����ѓ����l�_�O�y�OϨ2��KWA��D��k�l��-Ʉ�H3�bϳ�ѹfK�/�u���l������{����p�s4	�p����n��KaΔm��rŤ�673J�"�����u,�fPˢ�%�
\1���%HJ���7��Tay�'	����S�8�w<�u��%Q�ɱ���A�G�|݈/i��M����x$�W\��<D�wJ ��9Z(D8�a���z��� h�p�fl(N_z�wT�d��D�x��?��L�	�ŝ L�­V���os�_S]��W�B�݄P~��0��T�-S� 8K�g�����#W��=���:��#�1!�2sB����!�����v��(�B��q.r�����ax֭����f�Ép9����;�|�}�"��]��}��%P�>4�<>��1��Y��t���@�<mu
�H<~8�{�|�}�*�[O ��C�r�~�a29��=��s$'w��_�֑K֗�-l2IL���,��~���i@"�5���ʙk^[AU��p�/yĹO7�
���g�EQtv�gY��Z��ť�Ѱ
O��ps���1�w'����I�E��ה0��6N!-/�p�(蘇4�E��`�+&�DȈ޽A.�yrCf@�L]*F3J��kP�°�y�@ ����۰������ܘW���$��p��OsM���4��(a�W2A����U9;��R�s(��#��ׯ"�B#��oD��x�QO3��� ��z� JP������w?���[{(��/� Qp.sG�j�Zh|Cph�G�=��:�=-���8d�n����HG�c�� ,#��>z� :�F�����Cz��Bv;*;{�o�K�}�չP�t�w�,�@�a4ڪ�㑯J��b'η\@ѦH$�Y4>�ٌ�'��XQ�G_��M~}�T�(��M|!����O`iV>nH.�f��i�xl��:vǂ�w&�c�!�ۈ���G����(L�Bp܁�A/�m�.����ײ��x�TC(�}�;��mm������ä<�����S_z%W�>�e5$�ktid�3��lg}V�%b<5'!1��A,c1#b��T1SF��˲	�vԝ�6I�rq��Fܜ�������8��g	'�c�	J5�/F��(2RR!OJ�X�X�� 'SB�&VH�Đ���T	���:>�bZ��MNM2�g�ce�:L�m�[��uu����*4D����C�QL�=�G���FZ�-�=hoh���DW}BCN��!�#X׊ �#��[)�A���%x�����z�	Ӟ?Q�$"�W����p?jV�Bfcdg��joGRm��]��=���A��P�gAA�:ڄ��V|n����������*b�ƍ��x''�	e)�Ku:��u�Uә��'�Ҋ�ʘˊ1���~=Զ���� ai5�7mBJI9�rZQ�HR&D�W`B�C��$Ij��R�fQN���C��v�Rz��hd����)� ���Vw�$<���:APTD��i[%��2�����cI@�m��u�E*�g'�#M���Ol�`h�4�`㔅/Ő��
�a?ϴ��
�Z.[�����:u:qx��O�HIZ^�R���dȪ*!).�B!���I�KQv.2������JҰhV���LL,�Il�~�ǆ4�������O;G0H�0�t�,ǄՆ��aH'\�Cn� Lpx��B�.31�� eIZ�=�	��Pખ��"�N���63�e�X[�u�
�e-�M�K�����}��[�F�˃����I	���è��? x�w�o��C/@Ǘ���:0�Ǜx��A��'��Ȕ%]D H��d�3S�������A�YBl6�r$I���Tz��V�ÛY�����yp�b����А����G��~��*	�i�����T��PXl�o����B���M�Ҳ�(+��r�S�#h;|w�ec�iGi����j%�@�e�Q��mà̈́��>(��r�1IBm1��@L��2�,H�6]��._��U�m��dB��"�����tD&��O#�Q�?i�F
<$䶉Q"��t��z�w�7IbDY�3�� -���"t�6�s-�YPa���>�/�	���2#�)3��v���CC�?2<����2d��Jv� �_7�ֽQP-��`Y��eø��U���ē�H���x��y����L��s��&֞�����}�W~��� �+���_��>=��gM�]w�����b'Y��������<�4��"�!���Fdߺo�G	�da��:u���p�:�U�����[�K����Rm��2@f,LN{�xBP���+ �� ��$iL#�#�WV�p�Z>���ן�h�����dr1J�I#=-�Xe�c��F<}afl2���3Q����Q������^$���d|>��}�I�Iv*oG-Kܛ;C��N��t�b���C�\B�1�w��}'.�^�=,�b�p�C'̒�"����r��T( KR���5�	ݸ��"U+�v�j9��Ɖ\P����u�w?���Y]���JMn3�xg�&��]K%�>0n�����9���.�����z 7�S��[P�Ѷ��-.�W�bYN�Ga'�>�w�J�%r�3��]�[W� ��c<>�|�x`W45IX� ��O/��M��X��tzk0�jL#'�t�컓�t7�����s�]&�c�/���sHu;Q��Ǥ	�8T9��OI��VlA8��[0�b�8���	e���ain�����Q�����C�H�/���Tj��.����8��/�08�ga�r�tX��ŧ�z�L'����{f�{�zc�T��^�#T�x��YZ`@8GO �,ʄ�NN�� #>�	e��D\��C�|S��λ��ئB[с#,�ψ�q��e-a��k��_a�p��>L��u���!5x��(Ic[���;[�M����D	��6N!��$8�cy�0�_V8n��=�~��{,����=��b���5����+�������<���}�    IEND�B`�PK   �N�X��_8
  3
  /   images/57489f55-55cc-4ea4-8258-f1cf3d9c722d.png3
���PNG

   IHDR   d   .   �!�^   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  	�IDATx��\klW>3���?�vR�ql7M���aBih 	�F4��hS���H�

�U���u� ��[�(!IqS�R�j�4&�;i�:[�w׻���|wv���cg/�u�I��uw����{�w�4`H�b濙%�k
�ٟn�N�W�éR6���KCCC�v�����$I��$���|�aM�<p�@ʿ�Al@2vPq�	�L��᠎�jii���2ڲe�,��,��=�}��7�~�o�.>��~��Cs���\AY�)�1::J�XL�c+���b����0E�Q\n`6�?a�Z̜	[w�\��4�
�"���(JB��|>��}\��y���y�j�̝�h��t1 ��������X��rrr�6�������i��̏2�j����ee��UUUTQQ!���A�Xyyy
�(>ȧIp�bA� Q�������w�gQdvk޴��;�oN�G9��9c�ڲ��1��Ջ�x��^E�2�� vݫ���vH*�Y3J#
��Sv�y�F���|
!HT��By,�|�{�1J��i�D��O1ױuT�y|բ��j^ՈcwH�V���RJ��@.i'Iי ��L*H��ͤ�wyh��3�PN�������v�j�**b$}�O���#� 0ہ�����TZZJK�.�lc� �������137~��	�Ht٫ju��+�Q%���3�|��a[Hz�$������Vjnna�֭[iѢE��OD�@�c������������Gn�;�>�Z*�B�QP���u��r¯�����cتjz�p���OИ]�/3_3��_�����0��3�K7!ǝ�xvb4O`η�3��"��V|ְ�y1Q9n�O4M�.]ҷ
�"�"��0�M7� 1�a�$������h�8.o6j�0m�{�<y7P���'�lo&c��Y3���#�1����9,b �:Dzd���drG6� ��O7j��41NG"#�L��Z�4>:zs���H�̤�1�!e�?�>�|��b\�)��{|k����8v�#
`�:��ac.$a1�1Ě����2_$}�`��[�P
b��LwWf!�a	��T.m&� c�
��b��(�1TU�'��nJ#YɎ@" ����I�������@�������7m!�8�m�9XFB�|�]�{�r|����5 �h���T��)�!_���b!L��_YYI۶m�ˮ�>����0�}�k���N�ec>�l�J��'_M�ҫV]UN��������~����w���"d����.^�H�+J� 4���Lit��g�-[�M�����A!�����g�v�|����vwM�I�i��)~�9��(+$g]�k&��+W��,)�U!Z� �"����療��D6`%��� 񋵩��O~�܉?z��G���X ��$)\��˺�|�k �������^��h�����C�O0	h3�w�*w�o�N��p�7�Ap��W>L���p��OJ͗Y_t�|����Q޾ig��o�7=!����?�)z ���ڵ�x �or�Oix��a���YN'k�厰�dG؋��\�ѣGi͚5�v�Zۑ�b	�+ H�����-̳�=��)�03qc�AQT�V�Y# Az{{EZ�������S���&-A���I�:YǬa��|��i��	igS�l�1�Ng��|�t�YA,�Ę���Ux�՜G�W����kMY{� v��g?G��g��lG�$��q��MI&K����l�anX�g\%�*c>�\�<��,�F�)D9����R/��]���q�6� �q���"�W��3_���K��9tn��w�F����6�m�K�u-����`��XS�JЩ���1B�G��������n%w���HԈ����{TRT�R��DR�����yqu�0�G�%^�1k�9���+�]��z��8�̿zK,�~�oJ�EXz_گ���JJ�"�d��@�ŋu�m��wۘv�iqa }|q>�t�q?q��v?�_^�����>0Ԑb���Ⳑ�]�z5����e%Is QN2�3�ļ/Fr�S�_�i YEx�~���2��,c�,� �t�b�!�!������"�z��5Q"&Ǥ��b������ҵ@΀�,��&����s�GI�X�e�(��܈��+A��X�`d���&�dd�/�L{�rB��bx����DVbĳ�R��Ф��7���Q�$eOrр񢧵1,���/��%%%�����l�̉ �P��������K�:���6���Z@�c��.
��=Â��g���O/Y��������]�Q�E�\��46�]̇������6k0'Q�}
�Y�v�+W>��Y�h�U��7���\��� ^��z�ϝ:uj!��9s&�����d�?�`]�ḣ��k��(�ǌ�Qbd����-�Ik�S�l�C��%�KX���Й��%vO�g<���شc�aM�a�}�=�
�7    IEND�B`�PK   �N�X�E��    /   images/85bcb663-dfd0-4f8c-a6ae-bb35df534978.png��PNG

   IHDR   d   d   p�T   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  IDATx��]	�յ����Yg��ŀ��x~��|(�<�(1�xn#�Dy �A>%.Dq���q�� "����"�E���2��,�3�UU�9��t��:�ôL��tU�{��{�v��r��(8�����a�kІ�aP:v�RZj�m��Q�,���Z��p:�M�w3�Z]%���Gƌ��� �l�)��&8�=��< �@��u�N�c�@K�;Ū�|����@MWu��u/*����Ցb�0�}��4jC�Z����?B	��Wb���07���B��7���+�����ڋ��@��>��컡��㈖♡i�@��0���n����"��mY�/�7A�,�̽͐��O�6���nl��<4�����U�e���`�Z���t:2Zа
���m��a��d�-�L�١t�טKd��).\L�N؈��:4�_�g�M�\�JYi���Q
��H,Z��Q������W��vg���y�>{�SC���;i�N��Y@�Q��Bq��w$:���	E��;;����+�ό�'ܘ�F����V\�5��j�n�0qD�,�;����쟁4�OeqD������fG6n��������W>~R�/�m����b���.H�8��B�͍��,�Ɨ�v��e��P��͚,�Ɨ�v��e�p`ז�)/��6�<\.��yV�8$/�U��J�Eg��L~�����)�[a���xS1B���1茼�7��F�S�j5�[��R*���}��d`�����!	�O 4��BFꭉ�.z�n7g|C�L���ٵ�*Rp���&i�4(��p���V���todPM�� ��RU%۶Q�U��Ѐ�+�b,*�=�7Ȫa��Ū~}Q~�m�I���J6x���v8�|*̃��l�#d�\-k�4���������m�dN��h�Z�������~�Ba��$S鼏���y��<掝@U'(���@����zT(g�P�<�݈�ղ��H>?�f��8r�4��O'�*��+b��*�EB)v><&"���4u�P_$�"�+N9:y�u�)F�[S��5�B�PG��_���Q��|u�Mu��R"HF|�@�?x�l6κ�7W@��+Z�H[ lW������e��<K���������B�7Bɤ��*���nA�SO�t��0�ڋ����-�\�LFp�a1*LP��LU�zY����x�xk����w�G2 ���%[ �"�0n�
C�4����N����
��A�t�р.;�С�������v�қ'���YQ΄-�l�D92��<�Lj	���~5X7�/u��f�"���l�'�9���֡�n/�M�?�[��!#H/�`�D�q�5��z1�r�Q�8�����X�i0HM�LqzҦ�脵c���n��5a�&��̈́ڵ�#Γ2�l��(R:������P��<���\�F�@:�Im���������ǈ��|x?��������������U�76���;��7��e��0�Kzp*\��[����#��F�&̤�1
G��L�;|�O?#o�-��j�gOH�D�r���EL���q����A��C豾��+#R
$��`��4�m'	�_o�G�V7e�2���&؀��`oJ���r,���~͖�����ͥWȼn�.���*��C��ح����f	7۵��W'W�O"���r\����Y�Zϱ6ڇ��}]�T�I΂�׫Z���3Q�볋��Ѳ�C �(=RSg$Lڜ�r\��1ՆhY[ 9�O����W�e1�Li�T ;u�bX����K�Y6SN�v����Q�����!�1㽾��r\��Q����-0Q�mH����A�D9��)n�T�h'),QΠ��ˮ���j��)6BϚ(�;T
��v���h��!F��reFq֖���J 3��E���g�����3!�m�sCQ.�Ο����v�^�ps4�#��D9ώ�lB����!��(Wm�C"Q�w�G��fI)��$�8�Ł^��A�`���ftf-�1$��ΰ�	I�r�OϏ[�r�؃/�����!l����)�:E�J�Ψ��\(;FOg$$!��
�,-ER_5��@�*�ʹb�^/x=t?���o��s����		D�D��$U7Q�u?�mٗrM����	Q���a�����6Q�EH'�0Q�t�qU��31���،���.��)��D����i�;�2��c� YfXD��m�\��&�6Q��`�6Q��P4D9ED��a�(�r6���r'N�܉�(Wd��r'.l�\ѡ�T~>.�IRz�$�B;$�ɥ�(����X��a��kq�Y��b@�$��Ê?��O0q�]�]�y;>X��h�l���r�&��R�H0�@U'�{��(�Q����e�"Jk��c����7���>Y��W���t����-�#�I�?�-�mM�3�phw�ն�Y��c�A��8�s�&��%�C�֩p�7jmw!�>�k�����۔(G�Qi��y��05�xN�8���B7����e�H��ϥ?�(�r�T��w|Ȯ﹅ �����!�QE�~Z��>�ǐ��1x�/��rs�i�m	��Qv�����R�x�l�o4���9��(����NT��������(�"fX۶[Bi-�@�z�B��Ƹ��#���w�[k��{6B���L���K.���)��8g��I��@#O�QK7W��f��.���x�q�;�B���&��V!�\$^9�׷�=�>5Ɉd�F7��[�@ɸs�0�|��#�RR��{���I0��-�ɵ�	�'~���,��(�S���#�o�}�c/Y��vC���f�x�UfS���@�c��WZ/\��)48���b���c��V�e/��G�o��G�9�1���^�eD���}~>�L������+�θ��߲�9]$�픓���SO�i]�fw����w�b����=���1��f	g���^q����P��|y;gdV��1���<t���6��D9�%�]�2wd�yBk�/}�F�X�.���:5���:,_��[oÿx�L���'D���~vIs}.���,E�ԋ�{<�MD��Mi����8�s�3��L� �b"�q����w�w,
RjMW�]%�\����:��w߳�[Ƌ2���us�� �/\L:}-B�}�O'�r�"!%�����,J�b#ʱ��o�&�SW�!�|S������n�se��_�5�����VpK��߃+�X.x����L]%Q����;�B��@k��Ybp�,L,3���Qa0o�+�@���:�Gi���P��$p5�E��L���Ӕs�RQW���=�G�����0�
�/�2�}<�5_�$�����1<cS�� ~�^�0�)D��˯�-��p���,�*��L���X�g����a��RRIz�vSP��<\�D9I��h+�Sݨ-�Ђ�8��F�������'H����
������r|1�s��z��/��_���xR?M��#(�����%i�~/���$8ٕLc���P�ll� --�D�rz��r�(�}*ܣ.��_���%�3��!������_���]��v���R(j�����2y��d ȁ�����[5`�/|�r$���Q���R��$
G7O��٫"1Α�'!��_�y����KS�U�N��?g���~k&$u
�y,�숽�6%�q�������V���13!����tI������z~F���C)_ʒ�o&Q�4�����f��
���ڰ1��@mM�cg&G����%K�%�N�=�ogE�c�14����/Zl�7�'Ga��-Q��NeCՠ��#)t�d2�:���{�������������=vL��_��s'�-ۤ�8�VZ��-}�V��.��pPR���֭�(l��CD�m{����)̗�	����C��NY�b�cb�gϱ��;Qr��i�]FC�^:NrY�fsPƫy9>�=��{��M�u���8f��Fme�	H��'�94
��-@��X� ݴ{���u�#���j����gP}�&�-�Ӓ\UI��Uk�P�"���B���('�����!�_|)���K��ΰ��M�7Z�}�wx&Ma 76k�Ji��D�y�k��wט�i����I(NKO�3���f�6���Eף�m��'�,��*��|L�(WQ��#�a��ЙΓQ�v�W�@t�\:��^�5p�G	A �z_txĨ�w��j|�:�f�Ï�5���������Aߵ�^SQ� ��&�^�G��v��'�+�����`g��(�z<�g�*Z&7��[�����R���q6���ta�͞%v��
�9w�lFh�y뤈�f¨�#��ӡ����Y��*7�SP��_&^�p��c���f�Q/3���֤P;US'�ԡ̡�P�M�.�Z:&��p�Dp�|vO�L��y^��O֩�5n����i>L��v�?|?��5�)=�i*B��%kˉB�MeZ1��p]r*�+B�=�Px�˳BS�]X�lj�$�%E�Ms�t���c��ބ��5���0��( IH�Ѩ���|��{�%�:�EӃs�j�ZdΙ�04�R(�ïG���+W�*�5���E���$��ӌ�h�p��sS�1ÿ�f5Ů��}LZ�u濡���d����R��?���"�:���G�o��y$Ǝp�\��;g�)յ�,�C��\�</ћ���M�5WZu��tr�p���9e��2�z����)$^.P;v��c���������Qҧ�Ь�؍��� m7����'���ԥ�
�\�&���qٵqi�    IEND�B`�PK   �N�XN�v4	� m� /   images/91e5cd07-2a88-4b0d-9128-72e2f992e16c.png�{eT]�����ˠ��Kp	 �Cpw$�%H ��'��Kpwܝ�y��_{���9s���vUݺ%OU߉��*��F�  0d4  j  � ��B:��Bt�R��`�H�oT=w �P����S�^�����t���6s�X�Y�Z�[8;�譅�(ʼ��u�����.q6�n5&��h��H��tҠ��_���o_���ݰj�9�j`@LT_�Z��d���BX��%����T�^�O?�ڻ������;�^�t��#{{Thm�+��j���J;�?��G,d���)���'eH8����%cG��q,%5'��O�N-J��dj, 4��v8?Y#�0Ӎ��?�`.�V��z1�O�������{W�8�^����ap4/~b^���P��^���}��@��-:P��:{1��ΑW LQQ���Z?���U>�Z���N�1C�]ɅS7�HM�3���?�Y0��sZ�ۅ'� ���%,҄nl!���wD���`G�b+��O�~������)����,�J��z Rɻ$�-�TR�*Q8=g��?�Ѵ�Y iEH$#'Iz�oY����+�a8=��b0ҟ�B�T��}��;5ʻ�;$"�;W�P��$⛩�4�_g�,�� (7?�Ɣx0@b��awr��`��1hdb�Ծr����Cq�Ӿή*�Ä�݋�q����LR��\�v�Bo�`�z�̐��I,���F�4�!�����!�
@�p3O�ij���0.����ZeE"�X�%<|)�ؤ!�`3�2����a�ƈH?��¸�$�� ؈�H�QGjC�T�ژ�B�`̄y�#����vm&��"��[B��IL����g"����RhY-��C	�
�I�H�VAt2�w
�Z5����얜����e���!V�?���>4���>*$��H՚�n�	�RBx3N�K�#�u��_�u�a$����8�d D��1�J3 7I�*E�ưdB�������ʠ�DJ�~7�S���yj�d,�8#V��K����������,�cʪ�c��C�������b��Z�8]| d���f���g���sj�=�� ��x��!�&1�r�Ӕ�`�co����#��&�Q2G	��~��^klQ�0>�s�5d g�B=�d�H?�JsVP���/�ama��&��?X5]�(b�Y���ӣ@��w���'�.�7igi੅�)0��VK��E�i*W]�Tu;=�,����?��7q.N�;�.��ڴ�[P�B�6��[T����*.E��ہ-��'_sI4�Ҡ����:���=8R���	*�+��t�}�k���7b����{��>҉"�T>CG����WV�Z�����Qʈ��^�	�?��9�̫P/H�"��w�Z�S�;WT�x�6��:��I�R��E���� W�}�}�{�*К�ì{6\m��%k5'u�A�lK������l�	u��4�x�J�r��
e"
��ו�+)�3�+�֔�OhԠЏǻ��qF
.�^�TȦ<�dJj�_y�8=r�v��g�E���0�ۆSkJY���{��u_�#��H
߾��92��8���� R�b~�4u1p�iF����".pP��j���{�<���ٿ��Pu��,���t�ڰ)կ����ݵ̷��xv�լ)���;f��h�N�y��?���=E,��&&���;�"j2y�0R�H���)d�����m ؉����3�.� �U���ցm�l'�2y�1����&T�70vႝU_�X*�X��ˁܟ룽�����<׋y(a�Bᇇ��|�է�/�Vē�'�)�o��@i�_Gx�����I�UeO�Tl��	j��#��Q�TӃkw���G�C�#�X�ƛ9����2 j����J�xQ�eC� H�X�f����t��tPԯw�A�n�r�7}���R��uNOǈŜ.�{����U��	��z��잤�a;��ب	��2;�<�U���[�0�6CZ�zP ��$�;�k���1�����-��&}��ܢ�}2Bsh�쫠R㥭=�?��65$꧲
�Ɏ"|��b��{����|���M��^�$�0 q�$"��Yo�Mp�+�ڊ2�#⫩�+�>�����J��t+��)�W<!��K<^�>�ې���YO=����Q�%�rpb�Q\G�vË}il�
;͕`N����Ml���`Q�昷�;��O�S̯��O��R�>�}�Jwɑ��mq^���Z��o
~p�EI�DŢ7��M�������SI��C�2�YWT�N�I���#��
O�1 H4��\ԶP��@�^bG�A6~/h�N�K��'����"��Uo3�0��i�ZI9V~�9�(�<�Yk!fӁ�4B��e���%�jכ'>�4��?Hĉؓ��8�tˣw|�AbH*:�I��-FѴ�����M��.�����`�(S>��H���ϳ�� 3�m�j�=�r��.��fm9�B���!�+�nc�x��#�*����k�S�B�������ug�.U��?_�}$J���wB�`\��PL%���17���/���[�YS>n� 0^C2 hs��Vw���/l|���!��}#Vs�s�㐻W25��G���c��޷Y���LU��P�&�:����-|ԩX�z�Z��WM;W���*l��@;���Mc���x-s�������k�*��}��Y`}��� Mx3B�CU��_�:������N�%��WO^��b�*�z�oə�h�B�cNE��<���½׷N_�}�������ڑ�)^���L27oL��Bj�q��Ǒ�9��=(�}���s���=��D��	.<G����ׅ�!�8��t�v;ń2��Dc{C�-Q�g&#SN���Ō��_ -M
�㘑8]U����N�˳6���/E�`�G��f�eG�q���0C���g��2��JY�!>r�D�]
���~Ӷ�$x�H��C$c�pG%�]��� ��,��q���=5�f)a���1h*k^��G� >�s�bQ�E^��J����1�uYL�:�
���'��s�!�9q?j6\(�x}��c��"_�[C?i<=���)�v�e�Uhy�Q~�g��
]������F+9F�8�FƐ,�D��觬�B�.�1	�?O�y(�D��y�Y��"�P\��<�[s����c�U��ߙ�*Z?�H3R�C*Q�����-ȁ���*7�HN���^gA�또�s�����`U�D�mɩ�V�-����i
z�8G0�U�d��;�H���X�95��YE�*�y�Ħd�{|ej2}�� ��Nd��tw�"t�h7���"(�2�c�G��ɩMb�jj�t#a�G�����A&��!�Ԧ'�b�l(��E��4&2;��l�(>T靳�.N �+�F�����U�;��}�mv^�2�vd�Ϋ�%���N~���d��\��U���=�����3��]b^~?++�����3�1���8���
�i����d�H�K��Ѝgb���I �5���ҷ}+.�
&��!�25���Ք&Fa�7�0@�_����}�"Nl+�q���/��&qY���G�5�?(*�5fvD)TP�J�S�Ȉ��PW<R#>Y���W�l����<+V �BE����֜w��]�/؛.��ׂ��{�K�ޤ� EO8[+��Ӽ� �)+��4ro���T��`!��'��%�յ�::� cc�ٙ�M8��g��J�t-���k�ja]�~9:�k�W����t�+��$�]C�3��i�޹��F��=E5�Smi�?�ib�3����<ȯw|�����^�|�^D�7��[�]]j޻K	$Á�P��&(�MT��"�6r%O	�|ԯǳ'
�7-���;_���κ�9ME)zJ��������Zc�T�������7P�Lʀ�DyP	\�Hw2ny��S���J@��E(r�e��Wɾ�����s�R����E��36:duǩ�bĖ�*��~���i���}��;`''œ�§��Ξ���{�5���ɶ�%�Aj��K6��rባ����t��A�x��9��{�i�tCk���D�ٍ���a]��Q��_L3��|�wϥ��[Pp@�G�2
>�ʁE��F>�N�\Tzq�Ҋ� ���#`Ax��<)h��N`\���A�6���ċA���.	��-UȈ������ἐG=-�|xȤ��9�����-�q��[�?�~�!�v�;���;M����O-���Ѐ��3�HM=q�/{!c�� `���|�ү�*OK��0M�t���"*����_,�U/�������/�NM@�n��_g5�7Pi-,3�$�J��z�#r���H�#�'&l�ΰ��D�8U����2i,����V��{#8pB%���eq}�쉻�� k:PJ�Q�C\��𙦟�
���F�=cI��lv&�^��Ɍ��~�Նc���D��m����fWr�P�*�Ƅ�&�L�+��'U��¼�sB_�:`�ɯ	���S>���/Y��cG�vK�O� 8���>|Q~	�頳����p�� �.�k:	z	g �Wq��5r��k���?(�k���R����z�����=�bR3u�%H'v��~����]��'cd��;��֭��G,(y�����U������AVc�m��}�Y!�\�uL��P�b�;�Lyr��Q�"�T:u?��$`���^	�]T���WF�����1�[�����1����l<}<$�i�@2u����`��5��ù�p�\RII #��Xe��i\N���j�X�k?k�R���]���^�pa�x63 ��IYd��HI��&��!vy�o��֩����,�]1���K�}�������8����J���7����j�������u���+��u�$v	���F�eo����J��G+�9\��c��_*q��>����w
��S]f���٪|���(h8Q�D^�:������E�'�e �?�7�e	Pn���I*6�|s�W%�B4s����E<���Ĩp�S�w)��:��@5��솢���YPH2U$�&hh��;���k!tv|c���+�s�h�u��"�]+g��w�TQp��̔�=��k6�>ǡ�k,!�+TEWY �%�b�[/̀�������2&ȍX�*uY� �z-��K�h)6/Q��1���)��Kbldӡ6˟�@ַ��� /�IHۺP�gO��,���|���M�LQ;��7��� ��ޙ�-�x���o����V(Y���ܿ���S�)���i�D��}lY��*6���괷�Ľr���x����.��2S�]k<����G!�u:������AD�8S:"�Y��||�'��O���,$�Z�6C	��X�HD��)}!Hvʉ�5�@C�p��p{b�ň�H|�
��B�}AlJS»k/���^���_��#��}G]�&�6uN+�o~^��0��mQ���G%��[�ö�����r�~��C5�������ͪu��ֻ��%Ց�:�����J��UD}�06��=�[���EjɊ7O�]�F���?��u�-ř��k�V����s���I�<x)q�`"��{J����a.|%=:Ol34��+T
��zK��sN��<���2��g3��6�a��м��� �T�/��s���:}o�G�AE�cQ����o��i��i�`#���\�&W�=�h�/.��قIR@�Z���<�m�ݢ }����15�\�h&fk]�A�ۧ~'�ڑ�CKn[����H�x���� �Q�|�����S$�%�M���bgu~/�@*�3�&�rQZ���HL}�G.,>�g���栊LB�'%e�ԡ`+���X{�(�N�9"��U�~�3�W��?v���"wYz�dρ��w�BJ�̅_�&�7����k��pxMnй�9te^+����@��e��ȕ�o��M��\x|�iW�A�S�'���N-�B#Iq�+K���oY��WeL��OMD��\�<?�nu�>�)��y,�Τa�>w�t
:q��� ���6����!)���c���Q+�u%��p�-��̀��{��#]�p�iI���Ϋ�cR��b�6��ѩ��!��b���O+�b^��|ޭ�PP����*�B|�b��H�{>��}�S��.�Ć�^>O���m��`G1a��HĬy[�LAL�:��V��u% me��P��Tw)%AF�(,��`M 1��^�>�D���-ə��,]���ȩP�Y7���u���C�6�9��4B���>IƐE�v�;'H��2�.��+����j^���;cZ]�Łb�c�;�"��UT��G9������ij.T5�����'����j��k�98bu��o�"���ۮ��RLb@����Qv���,�$pCJ};x7�	6SN%�=�jw����$Z�h�t+��S�̇B/u�B�R�9��2��W9�t�t�.�TJx����)�6^�Q�;Z�i�%��͗e�m��1D��ߧ���ı���y	����#��px[I �� y������)$��4��8��-q�5�=fHz�z@�� �z;����#�ȫ�����jNF��K�I��7�)S�K�V��#���?�?�[����R>����g��9# g�'�~��_jZ;�V@1h�I7�?X��֧��H�Sr کh���*��"�Gb��\T
B���Pq����gek_��x�9�q���H<�iV^�~�_)�B�E�ANW�A�ːKU(N��Z�ﳂ�L
,�[5���P�Sr��N�Twʇ�[sq��D�λ��Ռ�0�����y^���Þ���4���T��U�h���w����>�{�[�c��W!@j�476�B��m�  �t�w�:�G�@B�&��TVXk�ͥr/��F�jВ�*�꩝>o�^�=PiN�cP�U^$�H��M����y������'8��ى��\k�W)�rw�~��+�(��K(ݸ�[��Ҫ��rYĄ�ԡ�&p��E���?άٝ�55��`�4=���O�hÞ���ϛ����лe?�K����/���M��,h�qB�w��5�oT��e�mq���8���k�j�`����BVU�3��e��e���C4�N8��&��p��+�Nd�Y���1��F�]�b��Q8g`}��lAx=,�AHng;Y>����G�Ga�5a��9jh֞�"���ڌ�bl�Es����rЮ�v�i��ٓ6�f��k�Qk�O҈���J'=�)8��Ԗ�.&n��y��&P�E����mc��]Z���x �~sc4���K�+0�LA�iz��Y��`|<���S^K��48�% �%���k,R�7&s�vx����)X
X��8��0D
�B�§���͈,ݒ��\P�T���R��I�`�U���i[`H"@=����S����}�q�=7�胵Fө�_�bo0kF�2���}u�ΘɁ~�G�B��6+��o�́sA�	.H� �|����"�k���;CRu�'�\��7G���
��#����Z�g~[��J�gyq6h��;�æ>�T}c��#�b��ێ�t��jɜ勷R�}���w��o��%s�`#�_�*J�u�>��us�P<[��#��X݄�Ћ��?��ce�G>vX&|A�1��-�!R��6,Pء��a8U�yY���ܡ�0ֈ�B3Ay��F�F�.ۣ�!����U�`��� 0`�W�Z� R�%ġ���孥8R�r���ͣ���E�����e�[4���؄~۰����/��]��f6�Nh��a���B<S�ݺ��z���w)�ЦgOսQ�!�hkN�ܨ����1�.���h�5���U�w4I-��7w}�(���sz����L�=!���r�Jf�å"xTe+^U�)�c��VcY��\O! �G�G�ZpDYY	��G�>�إD럜]�/���4�Z�\����UQa�i��_�F�B�Ǿ���$~FzXgв:����?�hU�J��#�`��YSk[�Ys���!�o�ꇻ��Џ{@T.)IU �|���g�~/��ij�Z@�iK� ��҅M��X�"M ��$&�o�O�1�8�*�܎��9% 1Fi��5Ź����qҹѻ �I���'��u<لc�- . �K��1I~Ħ.�A��?{�0�e�/��������qv�� H�4���v���Q��YHO�����`!Pe��'��st��^�^����GQ�����L�9Ro.��~�^�T@Ot���qrDـ�[6F&��j_ܜc�����P=l3�.���a���A�]E+�dN��޼�w�*�y��`�t�I"Y�v�W��Hhv��%�Ĳ�������-"�/ߡ{�A�b�%>Lfd�C|^f��]F��V�OB�/�U��,�:{L��k˂���W:@�7:���PÖ9�}�h<��@�6,u���F;M���[鈈d��H���m��Yq3��Ж jȣ�����+����ێ+�p�&�_�M[�(o����@G�=-�d�U�����*�pu����h��XV֦�4E���)���8ڮ���[.I�kdP��J��<�~b���k %x��{���v݅��\�~�(�\���;+�j�ix�;_�8o&���FK��� .3کB<�W�-һ�t� 6o�p1�i��޷�g��>�Fw�<\�>z�Z+G���s�|�|�e��Q�z�����{F�=����0m�B05�<�$���k��t�8����m[�%uY
l�$����J���� �u]B$i4Ch�E�1��]�_эCf�lcs�6�#\��%Ej�b���cQ��he(,�=��	�����1O37Ḻ��Yy|��wмE����V䤑�t��N0�a�J3?�������q8蓻֫��v\;��mE��0�H��?��-X{��
�����b�]@OB�����~���d�QLu�>X�f�����P���J~F��B-6��[��#]߳�1�oRl+|Y�o$�O�4��?
��J��������9�B�$���ʯ��V���F�Cɬh�4Pf�ϵ� ��D8�<�܄E{�;�k�]��e��d�A%`�=No�#ɉ��/6@#_��O]���4���(���F��Z0�Q��[ZwIss�d�O �)Ӿw��}bn1"�{vxwU��ŷ� (A_�i�#�m�������ӣ�ϲ'b���v�Iv�^N�ޘci@rM,�#n&s���6&w{'8a��{�Z*�/tAH%-q�,�h����϶�x���󚹯ߍ����#��=J��}Ύg³%F�zo'rC����U�d|$��V^�N����_��ZJ=��=�KlZ1�]r��?vtXc��OqYh1�e�:n��8�I���\Hi�.�{�9���[�NS<���w��o�ꮎ��Vۼ[3����R�?��\!�[8-bw�D����C���_���;huǼq������ro�C;F5��Ng���V�.|�"�D(\�ߧ�u���� H��y��1r<��Rֆ�]�֞��k�T�s�X�YRgU_ʡje�QX-� �4-#��u0J��+ɮC/(>�G�6a-4h˳F��o猙sՐ��ǒ9u�X'+&]�!��K%��~��},�m��"*�����c�·f*1u�ۭ�oo��}���yT��0"%�T�~�]��
��VTdÞ�(!@��k���1{�<��,��rY�5�=�
�V���l�U��"��E:����H���z绡1�w�N4ܵ��"�f��?���=�7�{6��*��D����VZI<U���i�s�W�3�c�ck���*�6]>�7!E?b�3ސ�d�lV���&x'�Y"�fQo��;W��۝�[<�em�y�&��/ʸ��'q��%���I���6���;������r�d����I3���^K��i^&�ԇ�o(�D�{Q~@e��W�*�	���)���D|����o��uQ�D.
��"��\ԁ��큮��[�1IA
���v�� :���<F�$�I�h���S�(��Y�M��Մ<��F,��\�g��ݒo��T.����w߄�LZ^U��5��c�w�
�DN�E��������A;Đ���>�����s��t��c�]q�>p�!aV�U`a0�b�v,�m:v�ٻ����軱W�������n���|�Z^�^���_�t�/���E��`��N��׎��؞_r��j���v�2?bŠ�D�u�� ѐDV�*a���!m�i���L�H��!�a3��/���ߓ�k�;(`W+ k���K��ETѿyv�����P��`���}+暘7<Ѩye�cS����P��*�$E���Cμ������\��ߙX��K+�*�0ȅ0C�s�V���'����J)f������4�՝~& J�جcILZ����6ɲ��H�Z�qD��4[�,�����Q:�iN�z�A�n�=�3e��4����m���?b=8�P�w���=Zl�E��$�ܮ��=��y=.5�/���6��b�J��#?ʀjN��ϳ�?���ęт3����ƨ��c�Ҳ��dL���HĜ��l�9Gۙs+*�8��a8Z��\8}�)�o�&`�r�R�	?n2�dWR�{�|Ya�Gr)|�Y>u��^��+YK�b,-���i�gRj<�{����]8���#�~�=� -��V�T�����8=3̴�.;��U:�;;�n�ii7%���Cд6�xʶ���m]���%T�]�����������b��":O�JV~/�^����=qЂн��	�Ш��olii;%�o�VVb��O���}n����=�Hcy��24ifap��B<���y��m��5/���v�5E�Egݾ�~��Ǔ���Ӣf�����{�&�Iz��N!T���0�|�${�Ϧ�w�`tŹ�pB�����4n�5��W�
C.2��r �s��Ɇ`0�JW�:rajo��E"���ÃR��B���=G���'Ku�ʋP�!s쳚8�J�P��>����Z{4�?6�[�{8V�����P�FVRTt�������y���5�ʲ�^1&HĞ���E}�-I�;,��A�S�%�P��U��v������M����d�D����%�	��k_�:{��TAoz�;�j�2 �����NB�w�O��lx2�Gd��1���b�A���H���]<Rw�>��#%|�����&O��D��|!f�ц���&gٸ扄f~�_�K�j������6Zy���:����̝Ij3�M�ojz|��b��6�P
�5c���a�}:�ڣ&��=qdiS��Ew'?�߅�>|�g"ͺ��n�Đ����U�� �ꚴk	�y���.]�^ň�������k��5t���(�ѝ2��4G�]�8xBa��2�7����<_Z|���ҍ1�;��u�n���}k��rU?�\�r�����ҍ�8<�/���7�7Z�M�G�$_3E�����N� A������hu���u�Z�K��̥fb�F�Qe��lk7�Y�7�[+!��u8����,�Wi�
i�h���Y~B�ţZ�F���N��@�}�/�o�րN-��aG��)��.ua���mRwҿ_��ϊSURrV�^�G�o�AB��~.���,J��vtk�ɛ�Ƿ�ht�ݦ�����ꕃ�c��6�H�M���\L ~�C�b����_C'C}ɤ:�W��TۺW�8�����A=k���#\��d�O�+9P��}�����?�{��D  I�iO0-�n/aX��׶~]>u�keo�H��B} ��ͳ4�Z��l��)@�5��.���I�M����
^,�q(��Bc���?�);�cOkQ1��x7��8W	5��/�&҅l�9|��:��?j�Ǧ[TpW"x��/}v��w)�����9��������썿Ͱ��qp�h���)!�="/ap�.5��GL��(�V�ty�O�{&�)J!ֆ��7=Y�V̧���MH���:��|A��0�+�vq�pM{O����Q�w��t	�]kr,��6�C��3c�ɑ˷�l=9e�㟔�}u�A��R�ѦZ�ˈ�[�_�#Օ��u��xw(�\,=::��m�h���)!qk<"�ی�/��.;�O�2ȏ���Y_�~U��~�}�ҹ j>�K��&�v���X�1�����w������g��J���������67�-�k��$)!y!c�?��7����9
�����]�����C�	j�����{
R/��]}�
�Y���K�^Y�y�5!��R)��A�*�����P�CH���g�T�,�&c��{t0L/D�r�(����<$Ѱ\���.��i���Ɋ��&!�8\��+�J��]9�˔�M "�=�a+����ԗ�u�h�I������8J~�����i3V���ÀM�F��S��FuA�L�x06Q����p	r�J�-�����Q0�%ay]��U`�?~arxPV��'V>َ��,p2FI$�y��dt]�T҂�	���7��� �!��P?Y�~Hs�	�.�{�ﰊ�wy��?#��3��Kc��|s#��#�����N~{.9���
.�H5X�|�f������ ���j0�#"�O������ó��vo_�q��p!�EB���ߓ�**j^�Pi+�Rffx1��%���I����n^#��}˝��O��"���!HܧI��r"��_����W���Q!�PRS�SW�Exxۯ�6�P���|�2��*�V�8ސ��-?�|_̶��o���OC�b�H�Љ�O��ϓ�5K��e#�#��;��!�7Ϫ��h�����zK��k.�&��*��U̾0�d��gƓ�[���%�j�7q��R�����Ó3����L� R?/Vh��kf���jL�Ui��L"�n��~�v!�j���0�.��e�����q��A�U�4@a���{R�E��D�۩���M!'�$�1�9N=����YVZej>��±��3�("�����+�����p~ޱ�r�`a�D6wV�e�D�IN6b�%��+*�������!+�9���n��
��$4pOfkr�n�m�Ld�zQ��$��q.b&�o�Mv���Ѩ��,�^�������q
�r�I��a���i������y�cG�ŏLt��˧���R��*�!b�G���	$�کO�^�u�1��Q��8Zݫ*F�z�Gp5��C����*��W_d�hӪ�F��8<�Ir�p[wf�:o`9�RI��$V��g����<){��i"~(ґ������Z_�����-�l��SH���7��Q&c륲Ȣ�Ai;q���W���{��oqp�T�]	��Ym)%�o�ӿ[�ZO��TB8�9o
C�\��zk^�7����y�@����٥R���/�F��u/��#��NA�N
eٲI�/Y�����d�
��B3�
��'�}7��p�~"Ih�1%.3`+���D� ��]٫���BXF�;�,;�,�����R�/�;��".�6"��ڊ���b�L���?�^66c��|��$o8�ҳ����^8"83�����,����i�o�q؇ڔ��}�|Φ���.�z:�ɽ_A�S��B�+T:�3��E�����8�M�[h�AJ A0�����}5�664��΂���xMZ+�X~���sQP�g�u[�X�=T��aE��_μ@v�I�g��Xi�F��� �#V�����^���ҷRDF7{�z���AF��˕�2-z��au\z��ӽ�6�����=�<�.�}d�fk��)�*�-��;�N��1�9�g��m3:����wHz�mE������!����O��yYu�B��˰�HV�ab'��J���6�T�5<?�Xv�_�(ZY�.x��<N�k��G&IPV?A��2eZ?�*�L��h��5
�V������"��͞3��p�� c.k�{x�l�H[�~���|�GPLY�P/
�H�/����b�!|!��Ps,'UF_I|G��q,�r�Q�.ʕG�UU�7�����`��u��^$U���BP�������K��9��p��1�:a� �j�=�@*e�;�R��˓��5i(���l]e��9B�cqC�$[�vy#7�U:��V�mM�n�D�"�h����#���ez�����	���7{����J�«����N��cG3Z��=���8�ș�����c���Vt��D���3�?�c�qج��-���MS�t�T��~Z��I&����$2L8K��p�7*6:3��:9~�k�X��3�꽹�$\�2�X�����ߐ=������57]��W�S���U��������6C�Aq|?�5�`t{��hF��=���v�dL�!���(��.�gg���J> �[A0ؔs�^�	j�vژ�pBz�[P�_/9-\l�ܲ�X���y�E0��0��.Ż�����~��y�����.�1������,p��8\�w��4Q$�f�U۹{��|��O�)�$�<L�&��q��̔�ԊM��'�!Cd� �w��H/��� -��b�H#�Hd5t$�zi�����Pχg~��w��=����y�vT�<{�35�eR�e~
m�;�Yp3��;m((���;9��~I�ϵiEyWW�%1Y�GU��1����@y+�H�@��CJ	�ȝ�F��3l_ө���EZ!��?����/��9��-�#��l%T�!fJ?v~^D��3��.���+:t�	魩�(�}���zU��p!)-ͯ��2	��] oALЍ��o�S3V�%'"�]�D���H��Y�>5iϝ���F��
�H𡸭�H�^�s�h���1��Z��_4�mN2���7x���@�E��E嬨�Z��� ��0stj���I�1�͖��?$c�|��j�l�	�;�I;%�P#z��gs>�n�D@�<A�h��G�C��q�ᇥ���ux���)*hԈ��춇G@�Nl�b�cԻ��_�a!t"Z)��������O��'rץXW��#]�{ߌ8 @ߠՄ�-�mr�Z<��X�YP��\�U��bBZ#-bFf)\���AQEųmGq�ⶒ*��H��Z;r����� �٣��:���r�b������6(�>��A>1�4Pb�`o�y��\kV�V�G�T�w#���Q��B#P�x.��q�Z�c���-Ex!�l�F��\w���⬩�8h�і�(u�J?���P��OO�F�c�)���r�̩���Ó�Lߥ�G?×L��S|�:��Յ��&�!o��hZ�V�r)����P��H�̙Or���{�
�
��8eq�U��b�?w�����y�vj�%�g���^���}O���]KKD�,�sW�� �ׂ/���z����kok�x��I���SD��iA�<	qmY���֋!��\Q��225t������O��m��"%���)���.rv����Ƅ-��#��ڹt�@9�~X����y�N{��O�Q˒*� ���[hd�Ŋ�|��~V]w~�A�}sϳ�!��ׂKP ��yfb%��\Î�ŝ렆V@[-,j�R����uŧ���C������4��YX [&�����	�=��z�@5l�c1���z�FC�n(�����i����[q>4�ޥ���ċ򿭷��uƺ�tїg�Qt.��\L#��%��U��'�}�G�����;�x��/��ݚ7����M����I�%��jG�&��5�֋���wBQp %"-�at���*���ɳ봭9��8R����y8��CcE'��85�]�����#��=��Wl�ŔY�^���I����`6?�o�lg1�����EEF��z��m�6�C�%�������_��RV�����*-�oo���>�l/z{�5�x�P�7�����o�ɴ~�������c6��＼�F������V�hi��-uh�&��Q�ه;����k���$6mK?�3�-T����� F�PJg���(Ǭ�ލ��yҘ����U?!e~"�cY�Tmv��g��06�����t;�&RN�6C�s�6�Kfj�I�Rs���#ىuh��6��P1
����K]{m��S���,��C�V�rNq#�<�Z����o�n����+����J�^���G����j����,���DObiC� �6�TU!~<2���zd�¥H~<��m�ڀv	�����^���Q,�dc{���|2cy'�������ש�~퐻<9����eqQ�67�i�=,�`5��И\T��V��������L���n�h������W���x9WսY�2���c�<�ϘlB���+�p?ft��6�#�D�����Ű���ҌZ$j�o�@,���ؚ[f��*~��d�a�f�H>b˨'�M}�.r����P7&0bl��l3�y�]����8B��4�1���p�6	�$�<����	���r�rs����~s�вhv�Fd>�������֧֭��}���Q�����6e�@t~`����L(����ؒ��5���bL�n�[{kQ���lf�n��ym�rp�֎f���\;99���(��l^ʞ���;�:��蟇�]J 𵻅^�AҚj��9T���8\�3�����'1Kj��J��	���&]�͂FQW����+�#ke���)��ogV&�B��th��c^!�����+��j� qww����N�����Awww���!����߿��p`�7����U�z�p�.�ۜ��x7%+B����T�K�������+)��(���^����n�b�w+n��=wmw��8}����bY^��!�YbI�o��3�������P� ��V{�Jj�v ל)pJa�nGQ��>��R�d<����,b(K�o����ܮ]	)��٥���.b�~w3��3]o���m��O��=f�WI+*�/���r>���$���"��N�d�"7�;vV�uŗ�z���a�V��=$��P�^B�?��Z�A��>P�Z7�+�Lϙ�8�;{����;�8�$�'`?���Q�_>�)��T�6k|���"S�kF���,<��Ltnĥ��4([C!}$�--�Vsxk��r�%�o;��ۃ��3Վ�i�n�1��&��'P�1�F��L��yfc���-N",.m^%v!�p�$f��F�}���kO7�(�+��YA�������k���S�e������]�Hiii������W..�PT0� ⮩�f�M8��� ���d���8x���)� %ā]�_�~�ӖQ�yv�[�BV��V���	M�-���o�x�D����lxPlu�����@JS��n�DPz�++H_���̙�M|}˫k2�}�D%����)�#�7I"�s'�;NF��)!�'K�IX=�/IB��م�Ӛ���QĂź���T���>p����.��K��( ��=���pmm-���Wc��C'D`l���G[�JT����Lh��7��/?�.|,�W�pF��`_ �D�>o�����0�4��M���#��7��zj�{�޵4%�)tdki�]�>�
���Er�d��:Ҥ�y��[Q[7T=�I��<^H�c���YC��8#�����,������"'�<Pj�B|V�~�Z��؛ӑM����F��x�8b;����P6��ï4v��H�V�y��Pa�---����u	!O��P����5-���I6X����-��yvV��e�!�QN9\�@��i�*Y�!|�QJ-����_���[�X�@T�T�`g�,^F�
,z���%FL�{}�=�W:��{s�l�d�r�a�n��تL<Ƽh�������#��b�����0H?��n]0y��eMt�i����7ڧљ���Ȥ�L~�3D��',�ۡ��n�k
��P���?<�W�6��iI����[Z���pp`�HΤ"�*+������P:[_)�& ����rx��%��￪����o�k��o�uF��PLMM�ă��h��tf+.��!���c�=N_^�ir&�����EH%��B>h�5��I0t�sA�=�u��DB�cB�qm.�/h�oũ�7��K���SsR}�^ę�U�c�Ѳ��А�u����uБ�����7u�V�������0Q bZ or- ����I2r9u5ҥ��sf���ë�����c	
���Y=�/^?4���F��]������F?5���j�U�����'��������tE��1!�K��J=t����M�eԯt��< �ZU�V�:��^$B�sև��L�[��@G�|E�|���/i��}�Η��_���*��JuA8x�T����(nN�/��y�S3\jX$Z ����e��i HD�V��Aa#��K�R���즥T���j�I��cj��sd�y?�&F���IJX_�'v�wU�W<�[rj�,KPLFl�i�a[{��j`H� �0�D+�X��n<�ʽ���"�d��k�O]y9��:���9�ȱ��n�v���T�r��_�x��_�����
�p��t�ܬ�d��<P�OQ�P5ăA5^yՈ�:�!ۇ���j��;p����{T���t���B߱�A��)�s�lo��r��Te�F ���b,h����r��Jħ����zT����:�� t��X��i#���&38�:ː�	�n�Eɐ=lp"�L�� �"��)4��=�����
c� ���A�6��[�1��m�����z�ֽ�{����.w�L���I��k���I5� M��T�������K|>I���d�	o�J���圁�c%C�Kio����y���N�����zF�W��Ӽ �!ˊ���8��<k0���<`����Q��ǖ5鉫R�D]����_!�s��[�8Ȝ/;������	<e���2��N�Jt�:a��V�&��+4��D������S�p�L!�έ�Ǽ�Z�G�Q�q�b^�0<.��2F������8na.�ta}nN9�,rwB���2�)J��5�g��Ks��كU/
Es;�q�k�4",�����%/9��ӗ�&�d�8�b��t��V��ݥ(_���{�K�B������j�,mP3�@��b��- 7KeFFщ��
Z�v�Ŝ��ضJ������!.�3�ʿ�iyԢb`g5� ������J��_�o�$E��L�׼"�[z�OUj�n����߫Ϙ�t"��I����%��;�Y�@u��KG�SOG�1ăVfNKF�SF��Կ�pȍ��Bf��Ahtn%Q��9���D
��R�:��X�]n������`$zm���|g����ؾ�q�K�̄��({��@�iY0F�$
��=�Zi3�qE�,L7���|7z���zј�f���c�znIL��3\F*�Z���9!#Z<n:n��9�9&〪9s��/I0�g.x�NȤx����*0e�b ޺�ĖT8�L��\A�ʈ�(�g0�������FA�Q�a	ѫ	�F���y�e����k<���ۨs����@]��㳻hA��$û��fdk���~���,����+S�R�4�:���M��ú"z02�q<�k�v�ʑ�H���U����p����iLI��Vj7�;���cI�bs7|5�?��*j�\j�ײ�T:�j��\͌L4̇�Q�N\������/��k�`;1�����4 �G�B�g"f����.@AVhͥs���r�=���G�?ت2����S�x"$���h<$��Os|��nQ�{ �x��Kg5�b��D�ڬД��xJׇ�1"M�C�ʬ_��]c�T���`�V\ōy����*B���9+�dqW��KR<�i������r]x4Uw��k��}�FNb��%�qt:6|*��P�{�O�s|�LP,�� FƉQ�La�y�&U-��u���@���Ȅ���p�n^]G��&{VZ02J�%�)(0Qc�:fb�ķ���@�i7V���3�u��q1��\zؾn�Q{\�T��b�Ϣ?P��8�܈#�D����˿�W�����u�tu�S�B�i%D�l����P~�Kt	�iRF� D�1�-):0|� dpa�a��w�U]W,l!�<���
��F�H2��U.��,�r7u���.I�c���,�pV�"G�ee0)0��GA��Da�|����Ad�%����r�dɄ3��p#�#㇀&��
o��1��[^���U
�f���c0�)�L�A�ą�de�(�ŉ5�~�CG�Gxf�Z�#��r�D���ķ�F�S�N��jG>f$S�WF�TP����a�_W4I�*�׻j:�yA������`�j� t�$F�1�Z��ʣ��x�����8M���g�M)e�e�sHR�Jit��cR�� h@����Kz�u%��+���� !�����b >��H��(�`-\D�b0*�(yT��1&������a�����.c��7���v,_4�"�����߽�ĉ0)'d�h��_������H����R���~��=�+��H��T�	��4�~DZ���3�F�����뿘��z��H����{%0�1Za�p�t_OЇr�>g"�[�6�K.�*���+�FNl����q���k(5��F.�豮%�0'��f��Β���&�C����G��p9g�`5̨�gnFR�	��(���;U&}>G����1h�	����tp�b��!2��3�v�x���G��ߡN?�P�-|�ߙhK@;� ��33��<6V<Q�#�_Q	�8QX2�e��%ѝ/V� X>�:�+����o�6h�Nk�=F�YnFt�AKC�i�J����ލ&��Z����rRG�x0��*Ng�ܛk����� <M��P~M@��+�\q0j]�jG\A��=HDv9l����-�m��i;ziZ&GT)�;n.*g۝�ߓ4�ɐ�(���D���	��D��|�E�o�"���C�՜"��)��NF��|�q�|3Q{�(��=�q,X��\�f�s#S���}�MW�	]�:�zO��ޜ�Z�����A4$j�%u��wPh���U�������J?�'�*XPvH�Z�H�̱Mw���L�V�� �&��F��K�*Z�x�j*T�o_ݥ?������cO��
?(т�^6ph���5B�W8"~ȬI�'P�<o��ʱ~3M��)���؃ �1۠|5M #�n�r1��k0B�W(�x]�χJ�Z�͟��p�v0t������� �}��H�Zi�����=H��=>�( �tQ�lCX�W^�����L�d�gb]R%��i���}��O�d��Wa
;����Z&���1/^)��kBD$�N����Iq��gߐ�ˢ:�{�=M����&���%%�����4���9޶M�(8YZ�Zb;�|1�9hfv�G,}���4�<i�ѐ����m~]��M�g�oĕ!^}^e�%Q��$��z�!Ѽ�&G��,��H���F�
K��ϻ�)s��HO_H�3~��c��bj��̛`�]��	Vz|
B�����t%b��詫Q�������ҏZ�b����g6ܒ@�i�=�I<$u��X	��v�R�6��Y��
S����%�O�Jԋ�
��g�/��|��]�/�g\m�I�Rc؟�YJԋ�@��!�؍;�E~���i��L!ar����,��x�o�7�E8r���<6">]��_�BS��&�	6�w����Q��]e�E���Ѩ�E��������� �H��������m1<����ƺ[���Ӥe�g��	�� Z�d���$2
�J���Ot ��NCTj%��,g {P�ɤ�Xs���Y��A��\����Ru �`����˕��/cGI�tE�f�TE��A8:��*Q6�y+�|����P�j�q@�\n7���P�J.v"�k����v�R�p�D�Q&���hMoQ.��fQ9�X�M)rتt$S"�n2��$��եwmSm�Q-)�^G㾌nl��4X l6�ئ�l]=�����rbS*�S���)�#���8���-�x�qkS��~vFj��t��(�fl�v�6�y,�b:���f00�X�,�k�XLţş@<6 KE�&��6E��hOe��z݅�	��̟���<MF���T�V�y��)�%�5$�����u��Q�k�D�	o&�����.=�p ��@��PIϞ
E�i�P�U?�&��2��S�U ��!����<�� O�q �Te�wlᖽ�ܙ�״���>0�u��g=��ns��BP��D�OB��|����<��*�@'��݉f"�A��t���+\�6��뤦LCm]M!ߐ(�35���2,�MT�������VL��?3������S�YI �G�_>�f�76� j�K�� �3�DW�L+a���C�q��,=$����_߻Q�Veqb"��k������n@o<��7e�$f���~�'��I�tN�	$��D���޾没��}r`��&�1tR($q����-*�����0(�G㏃�d�Q?$\���7X5Y���؇��fm!L�8	~�\��9V��Da~f�� L����ig�s����=���x� �84x8R��.�*�O'�OP��_M��HK���^u��x���x���L��X��1ߥϚ��$ܻ��wާ�ʧU�[]�T̎��j�G�u�z
�E��3v���9igeW����5����z=��������n$�X��N��8d�kqOqH�����m%�|,{F�������'�c���[�)n�]�Wm�Z·� FN!-_���X2�|pdCu�ob^��}�RfDy�>j� �JX5�\����*Q�Z��?��"�|��^ �:w�~�~�z�s�|D'Gf<剜i�����z�6�y[����6�"tw��p*�D8����y;E{��~'��ZC��̮Y׍�=C��U��ˢe'닮��ʯ����"��A���$� ��{~D��	Xr�8�L�\`�S�̎�c�؊�Gg��<̊����P� flL�jʹ���*��Oµa��+OȈ��T>=�±S���Ny�:��[��X����~�yC7><��{�h���:�2��26웈�Yk�x�W���l��j���N#v���=bܾ_1��wR���۟�S\k���||L��o��I���v�/���j�{ ����z>�,���D ���e'�v�G\8`k+�(�P��'��h0�W�+̤�j�*�qêSu�h�cu13*�D:�N'Z��!���A��E`���O�5C%���Ꟙ�{�z���Y&���P����?���wF=�o[n��7Y�p5ԓ�U���`��b�_F�U[�`��3ǩ<M��f8��](��c2r@t �0����.N��X_��_�Î�*����Nn��ȇX�ݜ��Y�������&�P�S��u;���s�I�k ,8ks)j���������}� i�~#o�g��~�4��]{=�*�Ki� �!8����=�1b��}�1Sg�2U+P2��L�˿C�5��`vu��� Zv8"T[�r%qW˝�D5L���D'�4�~6�,<T%�\D^^�h��o�1��#)w&�*jl#}%�����rp�XA������O^>�����y��ŤL�e�B���#}����2�=�}<��eḦp����A�Їf?\թC��0���4��3�-zN�o�Xy���rw��e��D�нM�#w����{m���_%�I��%���j5�}��)�9���6abT���vD'�i%A��0��k%}�wT��Ɗ͉���W� ���)dF������4�t��� W�0�=�Jj�\�,-G�Կ�Z	~�2�Q���P�P�iX$̧5�E$�8�b�R��1�7eh\r�+�!g���}�8�429x\˦�x[~�E��I�ؾ�g��8��`�������ha^7bFvqI��;:�0���N�lޱ^�o��?Еh(R��L��ȫ35C�t{�����I��+I�0zu9qII�²�-�e��fh1��H��`֩�d,�����_m��((ŵ�|p��ߙǧ��� ����Vx���[�����	[��b�������+W��ܨba)��A[�^�۸8�Z�"�������Xm��*B}�3Rb���y��z!N�B����%�)ma$��Cp���8g�\��(����'Vk���R	��k��R�y|��#(�$j4�Z�_�N�9)}}�;�+�#;��y(�Z�7`�%~�m�4y�Q�ɳ:K��\(��ݳ��!�H�6�}�ǚ��X`����.�G��1����׻ƒM��	��0!5?Tt$/7�eև2ɋ+jTd&&�y�ާ���5�gw�h{`�݅�\m�l@�T�:����Z�U�HIea���3;�M"����tеƏՌkQ��L�0*��1�6�"+q5H,�	f��ě��:7h��iE��η4;'���\���C`m<���T��%35gx�h�B<�d�P�i�lm�\�y�� KI��Et咿P�"A���l�2�t�����im9�J�`��6�߈y'_ڹS0@�-���7QRhԻP�\^د^�v�f"�>�a$u��-�	�[�[9G=���Z�=a��Ɏ���L�2���C�ZX�G�`�	���@�1���Y�K���S���������t�.���2�8FM��N��g�#�5^.��ِH���S0�*�ϯD��N�H2��ޯ&y����q��z�]%���򢍮�M<�Se����YJ
�;���
���V���g�k�1���_w9o#����߶"�>�/Mt��$�	q��F�|`�W<Y���s�34\��7���6��]���W�Xъ������HH�^�*5��C�ܭ�2���	iB~7m��N�Y�$��E��j��so�P"j܇�K�Z��ԩ���̣�`3gy�ܶK��� �� �ъ�6��g+0���o���t���'> 7�c��Su�����:��CƯ�������_�}V_���Hv�Db�䇪�lu9+�lXN>ZyE"Q�|�$6P��HBl� .���bwN�Xj�'	}���Fo>�]�:�/1qM�Bc�1=AX����l�~��
��N��wu��e�b�ԏ"e�}��n�,�5�� n��b���nwt*�(2���e��/ԅ�
�f��)�i�;�{�60�·��[+��?<6F?���o�~�ɫw2���޵�A�)KA���e��S��_R.#p��6���` �'?Iۦ}�.3�'�;!�"i��_��;�/fq����9E'ey�d�Fr��!�e�S_�D��@�����zW�ER�{>�).)u���u�B�*��w�������[?�����6;ﾛ	�o�����&s��>I��(�M��B��A��~M<D�↦�bq�W$�N�������<�j��M?��,�m����|\��G�OV'ey�[v&�p!$�r8��5�0g�����䣫�����L�P��cl��nv�;���}B��p'h5��C���ˊ@���R�j��O�|4���Z��xL��xx����^�t���.�`3Z��IȦ�.rsRI(
σQ���ri��;����1KfH5�uFEB2�̠w#:4xg����Y|��fJ'�j����&�h�����e�.T���D�.2�x���a�u�%q������fH���D�G��\�'�#�� ���+�+׻���_v-B�Eļ����k�[]v_���9���-��m�*Óf�׳�%��K��Z��ݰoy&�N S�n2g���<R�/4�]['��v:�q#`�?��L�*؎<	����V?hs�4%z{��t���}����eQ����)�;O�>�zbR[O+Ҫi��3=�9z�u?J��d-�AR�W+�,<ؖ����9Ӱ'���Q�Y��9�b��?Y���
��	�'��Đy��Y�v}�X��',b��o�x��p]��	�O��X�ҟQZ-y����<ʵycxU�T(@A�0h)�����0�@yh-[����%D3�V�r���3HP���S��ŷE��#��FtϾ�;!L*,��m&U�i;� +�B<� /��H?�l�`�Y�K����p��8�=���v�Z
�b��mt�&��O��Y���r���]?�1��o�w���l��ؐp����L��V`��d��%餓�&�������T?.$�z�F0C��e�by��p��$���F_�X%ϙ�����������	�?5���ml�z�������xU��~�������ȼ��u����g�����ޥ
�,f����jsU"o}�LGٓ}�^�X�P�x���hM�0�4B �cS1��o�s���ݐ��sd%��Yzl�ģ���9�*`�kj�kNU9<]	�u}��o��B=�+>z�Fr��_l0�v� ,�y]�?�Ѷ�wm��-!쌡Y��[����3��������B���t3�K7���#�� !-ºK!�#8�s�*���Jp�ۗ��dO�a[��[���" ������ǄşC�yQ
��<#������X�����I9-�ܘ+��Ȇ.Wz������D��H�N�7HZDW-QK0�.̊O>ϻ���Pt�Ȑ��B\6z�՘�D|po	�X�'J)Ϭ��1�svTӣV腀~��K���S�NB�83q�zJ�ז��گ�á��r�o�Q���hͧ�|&��0@��S�j���|�{�\'���Y� _9�B�O�P����+���[Ԟ��gš�u��BT}_� �J��A���O�X/��)�p
X��% ݂�	�� �B��
ε�8�s�gF�I"�S�j�w��j�q��?�E�(7kOO�1�m��`m-���K��<=�ѣ�t,��8��?n�zQ�Zʙq�ˌx��A��z���=�E�H� r�[�(t�7��V��K�M_��P��(��ة ��c���x����$L!�D�j/������#��'!킣]�]R0��^9H�*l���ӽ(�F%��'�:��֭�Rf�C�r���4@F�S�_>>��BtU��t�s�Dwe�ި%�������T�!	�d�3sm	���(z�?�G���R����z?X>��0E����6��7����C[�;0��u�����=����Pb2�����1e;> x���p՝��Ƚ1f�q%��p����'ȫ��b'�J��	�>F$/�Fm���P�ˑq�_����HQ�A�i��V.�]�-?�*�r���Q5�����a���c�K v��^��~DS#;�/��(��~�����Ϝ���&e������\��R���݋����^�z����jOvS�F�]h��-a*/��T�J�eFc
N���~/ˑ~�Z%�s1�L��/(R�í���н��Q\���ҝ�u�uT��ܷ P�;1�=|��5�U�L2b��{L��$������!.9���!+(���Z�R�� N�-��S�`�[���^N�;L,8S�\X��s��0�JG#(t��ޜ��ޗ0C��O��$<���\]5u!��i��=)%��L�͹�:��z�t6w(lW�b�Yn{52�L�f�4����
�.�8�ղ;��g �:f�d���r�m�o�V�ݜ�'�	����:���6_�\i
�����b]p�~
 ���;j��,.�������f�S��b�\u��:����Nl}��[��tE��jČ�{/�f8��)b��EA&���@ļT6�axXퟔ6� aRvgjtV�H&�+�K3o;!��Nkz�1����Tk����oN�P����7���uIl�,����̮�i8{z��K�'�U��y�/����,|E7z������zp"�?��z�U���k���|֞wBp�23y��� ɶF�2�(x�N�[�@B��LM�-�K����4!2�����e�h�W����G{پ2�ha\kĎ_T�Mힻ���d�X�7t$�́�__�c�rÚ��P����ƀ7��Yϓ��y�0|�> ��a -�s_��ȭ��b]݂S葩��|81B��C�5����֤:>�K��,GR;>�6/d'�E���(�|�T���^7���{:+����L}�i�.���ʟ̸VF����{�"��v	��_]�z�~K��Z�){ի+Q��'A||���l�/�2�D�9��'H�;��;���`4q������p.���$:V�ʫ.�� ԝ=�pei����i3�m�L���JHAǞ��K~�ֻ� �����,��T4OD�N"ʹ*V���5q��/z2�+�����TO��D����}F
6�I���/������l��p�D�4W�Xѳw�{V0t�|�E3 ��ٺ��]�D�<��g7�I�(V2|�z�[���m���M� FӼ�д\�]�}%5�N��ams����֓��?����r�E���k�#x^�<�5����
ѧ�4�"8��^u�l�����4]H�$.��Y�?�ŌUNT�r�IEq����Y���}�n k�<�����^�W	�w��ED"x��-��ʬ�����K���ZV1oj�0=;�{�����Qz�͚R�c%�ps��VX��5��L�W��L�i��������D�rP�R�3��&��]&|������b�HQML�0#Em�p�zԩ)���Д&m�Ek��B�)V$Sv|7��iҸ԰]i٨�aI���p�D�&0J;��>�P�ɂ?wo`�-��?��|���?O>��R�y���>#���L|�Q�D+���ei���.^$t{��&.S�֛b�;A��`��#YƷc���A\�8���7njp`O��ֻ���9�H�]�O-*ϯ�a�Ajj�#b��������@i�۰R�`�Ǫ�i��˭Xy��
��@D禉c�1C�ޘ�m�+��[� �ǫ���CTw�x?���i�AK�~*��02�3����T�Ԍf͡}��tz]&��ސ �h�n�}�J=8�;-mF& Rc���B�H@<�1�,uGS�O�c�E� �6��Ƌ�tN4��{�.Q``��z�iP�Tfjڮg��JKd�ع���u^.�t;�y2����4��e�A�u\/������3a3a@�I�b��V��Q�2�=�{���������f�>����`��[~s%�[�,�//0���V��~X�8X�v"|�a�*ணf��_��6�	Z�HZdqrO�?�n�-�I�w��6�/u��!�6�j��е�	�J{ �q=-�L�B��t�W��;n#��f�y�rÿ���ĿR�T��v�ۮm��O��=)�R�PN^�������f����z-��nC���B^��0���#����Ķ	e������שW�j�e�uX$�[�s�ß�S'��g� ����<��02e߇_��/��YA�HA���b�
� ��O+=����LȞ��-52`�T,n٭f�_tb$��!���}~�����l�LQ���9y��݆fDp� �]:?��}M���Ǒ`1�^[5���\P�bu��Aч��A,�s��7�#N�7G���52|7��<=}S��i4(�D�K]F�\����9�=���YyT�<~)��ft�>�ּ�,0J��y�Zp���@��.��ΉgS��R���:&��C��+���`���"d��*��d`C�'�]\��}`P`���� ��*NA��hj����E܊���ٓ���@
�nm��J��%s�Au&�%WD��3��Z������BB�{��V|H���i[8z�k�	#���w}��]ZW�b��G:�Bݭ�R%��������JB2֑P��~E���P9������\�d�������E�b��)���g;Wq2���6�=$-5��w+^O��R�%�Oi�^��$ϕF�y����:D?Vi@h�bi��o�P"���t��� �n��=9�{�d6fZ������i�o}cԦZ��~@��\��v�����#�%,��x��Ɵ�����9S�O����`�aV�O�tBw���y��Ƞ(q��"����"O"�?�[�p�p�RF��gC3`f��#��F,O�K%4pp�>��y1�)8��
����+��o���غ���8Ko�8V����}�r �J��L��,>3W��Fd�K�E��Mf�Q�R���١��nt���E�"p:(�-9�Rb�M��h,qU�$F����_����%��"��[ӽ�����4k�ղ��%g4Ӓ�tp�Dj�rs��	�aT��T��'4m1����`�+�48c<?���2��`f4#B��kJwhnw�X�[M�!�fsԃv9�k	�ԂA���EV���[=�:���Aiɨ�TdA�N*b!�~
�:�Zu�H�b@���=dZ�EJJ��YDƀ������ᚷ�s��!�g���[w,�f�D*����qU*E7�cAi�����4�=���������Ax��uw�4 &�^�'�Q��]Niu�ƈd\��NS��ɀfo��*��?Z�T��]�r8�OlW�f��̬�_�ޜ7�fP�c��ҧ|^5�?Z��(ˇe`	Nu}�cp�`A�V���7v�ӑ��yi.r��b�\9n'�AV�j�-�\1�n\���J�"�
e��?�����ÿ��#S�)��kdWb"�c�i1��d܄E����.r06��feܯR��V�ǯ�k�����W֥��L�î�[j`����#˘��HJ�����������=!�'��w��5ր� d��׹����U-�&M��\��=P\_�9zijf�-�{��U���(�Ug�mX�v�s�)���q!u��	�l�p�߳uW�8��� J9��ND{I�=���BhJh%�j�m2{�~\�5(rzӎ���PfG�њ/�W{��/@��0$��q�!��n�͞5���CyƏI�������na֤��P��_N`C����=�U01Ћھٮ���ô
��f$�:��P�k��I��Vg��7���E�dQ0����[)�y�z9�A�v�$�j�w���Ǉ�&r�+#����V�G?����'�B)���OQq:�LBr�E}������`K`��1��z<��HPe#����Պ���Qr��g���8x�x�[�Y�4�d�E�`��.���L�c�����ّQ�d7�jN�CL�	)����e������kM#�^@���J,��K���o0�e����wEy ����}�q�������iI�|��h�������2�(�����6O{-@T3q����7��۷yu#~��j�,`4�Y;�m	�cϷ�v�Bm��8���%��%�A���qo������B�@P����vs�B���h.��@�ˎ3�=`)Ӄ�;x�lk��QɅ�OK��I�/����n^L�����ӵ(�ʝ�b�V�*(6n�q��bb"�W08�ޙ�>n�zj��N62����f0_��A���UE���r��W?��y��v��{&}�`b�Y���b.���,����9p�(� q��~�jdl����o�b��BX�1�OE����Y��v���?��Kٷ��P�b��&(&U=��)u_�_��6h�]���4ႀܾ�U�:$�G{���GYNK�q�j��CP�����X��!�k�_�p��"&�N�*����9�n�#�G nq@=��J+x^�$�<8����SD�x�ޝ��@E���0��e͞�v�ev�<�i��ܫ��|��kb��T���xn���^9�Z�����7󀨟D���d�w�Z���\H�US�4곁�!JbC��[z��^7o�;�{�旞O����}��|�<���3Ç��a�P��fo��a1���c��6ҹ޿#�C�,Ȫp���A���h��.��J'G��)B�S
<\nj�¹��k%j�.s��4��5�}�,Ȝ�B���t�F��"?�0�vW?Nf_I�?��m	:�7aU�z)����thI���\7�޾�T��׋��
?��V7�$�z����ɭ�觊�����
}�S������4P�H��+�o^-w��D�!�Q��V��Pߺ�>@�⺖����s�ϰ�e�g�%��'����=�j�ζg��fďsˉzW Y*��1�>$f Dx��{�q᎘�
s�FKk��a�B�F�aO	�G���n���F��>���0gEx\�;�����]���i�[6ˠK�4��8���;H"���~���MP�%OH����M�Cf��o� ��s6��yq&�j�T歫[��^��A�3�KSS�^׆�HgӨ�4ԃl<���y�Gfmχ�=H���&� ��2j���A�X���z+(��͇<�èb�)x=bth��$R]��# io����m*3I����0�NPz�>=��4D{��3���(g��`���!�Q'G��5�W�_��|��	%Q�#���5�n��D��R㮪�t��-E�W��?�M7�C3> �Bn�
Oy�U\�9�ָ�L�Ń�jm�b��)D��.LT���Ί�=G�A!��'f�#�O^��Ԥ������7zҸ����+Ϻ���r��-�Y�"zk�z}>�5�a��3����뤔F/B8*��!�2�H��u�@�iOd6��Տ��߾�MN9
�+?�etJ��4���;��w�/�J$b|�׏:m�C���MyX+_�鮳�-�B��7w��	�J`��\���uw�Q��(�-߷�ک�+n���G�]Q�� �����
�9Tɑ���YY�^kKѸ!��i������6�'R~�
�Vb~��:��fAD �<z|(�z����T�	-���๦��Q��}L�of���T��fmgm��b���3�G�`8.,�=��ż���쳿� ��rŤS]��D&}>�϶�ܗk�R�k���Ee�{�,���Wv����[�6��U��:��wu.ln̯��-�>f�8���^�ػ9z��pJ��Sz��ݍ� ��	<�.����'�Q�����j�E�J�v&ɥmw�A�ef(0FB!�ڜ������u�m��mz��Dڴ)�3�������~s6(��b�*Zp�,�v�3� 6�``���$`���Da�d�2>z��?K�������dI�e�\!&�vʵ~<���3\Àh��t����)���oO��*⎬nO��z}���$��=�]�z8�OU��)�Nأus�!��
:	�=8���u����)����\��`��<��1��r��4R��Z�{����W ��4�^ �������!������	��w�<��v�|�{�
�����鞖sfzz�	�|w�mw�.��wZ=6�� �ջ��h�<r�x�D<n�͸��^�����\����=C&�vs�rȲ�#�[��߫�X�����u�.X�a}<�h(�/�	+%�q��F�֖1�U����	ފ��!T�\I����.`'D�ڶV�s�3��y��i!*���DL�B�#շy��������1d�M/�$�4�8l�{��&O�f�RR��{�z��wf����'�n��k�����������{j�9їӎZI}�S�˳[M������q5E5K�:�A
��sdwǪ_ie%+�W��0�5�"F*믖��և�H���s����_��-�8ǜ�~��`c+@��7��x������B���Z�8�m���j	�wv�q�!�� ���æY����|�1@dc���$�G��t�B�{PCSPɏw���4�BJ��C��җw��r�Ը>�5F�㺫V^>�G�6lY�l��@M�?D��kえ���>:�/I���Y����pp�K&�����w���0̍[We밚��:𮦗���.Α�\�v�� �TZnY �#�]�&eL����H�A���x�x�y��N[��h'�E��V�Zb���-D����|���x��	���\I:Ǚ3��SC��h]u�%�^3�n�u����#A�Y-G¯�s�����Z݁�����5�ߔ C7���$�~�C��!`�42�o<�!�Dvmr�dXP���y+���:��O��RT�Џ��hh5��x�VeKh!߶�o8Hi�Aꕘ�n��.�qfK��K��^��d]�Jt���`;��AO_9�e7M�4�s�Q@&�׽�L���7^��1J����:����%8^ RS��������{a/������W~����#��6���&M���mY۽|ޓF��I��E8���^�e�e���#x����ߴ]}ᐩ��
��#ף�������N�x���0��C�o���!A�M
�m ���]����>u�?:��zD��q�� ��֯]$
�������������ý/�P#�0֜�l���yno��q�8�GE�E1bE���K�D�5u^؈����9I.����P�D�����A�}:�Q�<~��8��l���k����k��J�if6*�Y3���>H�JZL�#kc�������R�F8�0��$]]]u˧@��i~��=w��x2�̃{�K��wM�9�^m�����.��]�y�/犞"}�̍�v4)�"
��.S5�˔O-�&ժ0ҥ5%o4	��9V�CYhw��KC>�Ee�gc΢5N[}���=q,Z�z`"��h:�
�J�ݽ�ܽ&8���:�`#~>ݎ>RQ^�C�A�ʿ��ڬ���5�o�E���fg^caipL�:�7'�Vwvv
h���n9�ӕ������<�~y��4>az
0S�pRo���(�/)�b����m��I�0�L����5T+H��z�>VĚ�$-��kXdו��!rm�T9bZ�������? �{S����+�l}� �tP��Aj�d$�sa̕�&5Q�3�&鶵��3b��|�죘�jS]�7���9eH�,t_��ٷ�J͛[r�QD�����C�lXp(�w񉉉����;��zY���!?��OQn�A%�
��YY��3���dd'�F�괫eddP}	��f�����Dx�C�l_�޴[��b_�2�@�3+A���YCz�?�X�.k�G�?&Y��`D�؟�L���+nٱ*J]�����q��١B6s�/MT�Q]�I��*D��"|e)��%�#�r�WQ;rC-,[؊j��a�<7wwwS�Y�OxH�E��E�$]D�?�c�>L��V��oʗsF��L���zvnH�W�"r���@���<lדwu��/:�����J�ێ	�q����*�^ ��;�+8��/k�̓�j��Rr�]V�$z?��qD�uB)�<?�d� �^SZ��A	'Dnjl݃�ˋJln+"Ȑ+�4c�P6[*#�kf[�q��j��9ǽ�#�$�N��0�*��vP��x�6AH� 9K�	�ώd��xˀ�'�O��,�Hn�~�p:�9dn)7����5��_�2>i����\�d������<����o�7��9@�y���f�T�<VS�8�By�rP��d��ረ�o�UPQ3��B�a�0���͔+�p�ڎ<��+i��zA�YdA-�-ftH���&�*O���T�˖�7�d��O��GJ]��5wx�ЮI�.}�B��Wuy�^81o7|LT��D��ϼ�l�^'ދK�d�`��X�� ��)cy�,��"f��IL�֥�xgAo+�2Ej����[}K�3����T,���W��T���c届�vc(�	���(�햙MS�K9�廻@���~.2c)�����=K>t�>`�q'�d��O���.C��H*OeZ9�>Am�}�y�{X�"Չ�������uC�廂wN*m�JN8@~��X��bE�$�����a�%�
%[t�0 �(@�ӫ�5�U@7�
T�|z_��/��rY�1	1�kq���}�7����������R������ɘ�t3#���٢���ྍ��MT��:�^�a�:�2��"�ܞWu�7��/�3/;h��a��|9�טL��k�$��ׄ�j�R��G��c�~
v��L�Y�t�p�Ƹ�E�۷<} 9��{-���]�L�A���N�d��++�`g�h���X��#�t쵼��du�.P�� �xb�`�S��H�%;�&H�<,��Tds~G�#D�bF��v��ho�R��}�@m''��'��?<� �#�+X%Xg��r�(?;���ճr���jw�V�²O�q�w�MTE˂?UG�(�"h�.��[�����;�N0!}�J�G�,1/��^AbІ���˿�8���a��e�FY�3���;���܃���J��s\�����v|{����n�(-�1x/��V7�l���
��?��@��}��7�����M]Zk�[I{���x/��KvT_s�	���O�1>S��9�*=Ls��>Ϟ��[�EO���_(�v���#�2q�/��}Eh���Po�N��ozJ�+�(|~?%���'�c���~�g�V�o�9�:���#w���O����-�"��sB�5M�j����G�b��w�`"L����[ȶ]5���.Zs�'F���ԅA"5�zUhuϧ��;ᬿեA�9`�ć	-�Ԇ�l��1���.�5�Րy����삭��������L�B )N�7���Wo.e��^���)'=�h�D�k4��s»�c.h-�����ףc���h�H�l�#
��
�~=���1ӈ�_��-N.�zD�7��It����t�cQ�
 �$!eE���:��B��bcʈ�nM�(n �$
��uZ���l^;`�2�{�wez;`>�����]�F~+��_�*E�r^�xF/���\;lx�N�G7�7���I�ȸ���%�U����C��pe��KC��G��3��?
L6�#=�ʶ!������:bh�?��F�	0?gZ>{ĵ�ckK�g�c]",�l~ $��Y�wl�ԾX<�vh߮��5���dh��0A���MS�L\I���׵?R ��&-9@���3�Ƕ5aXvN3՚P?���~/�2/�]���̟�މ��.ӴQ?�v/���H��/GyԌ�r>��VjZ�%��}&����y���X�-|�x���I~��,��mЕI���g6xHxq�a�<Ȋe��n+������1^[�떵���b[k��a #d�����3ɪ�d��X�+灟�,��]�GO�j���\��/8O:���Ž��l��$�r�_)�:����A��>����>oTOM3�Ŷճ`�Xc^m�Uk0=۽9=[)I���w2��a\�O�C?�Cn##��_��c �U�V��Ύ��E�ыv^͏�F��0hq�}��
q�:>��:��,��L��(�^u�[�P�(B`�GW�"��D�7�v�f8�#$F����h��߶	�
jT+
�i����<;V�t�r��ʵ&��y��+��R�|�3����m�3��k6���L�%�C��������T����3&�}��A �7�N�;�8�hԓ�i�P=K��S���?�4����Lc���'D�V���N=���~��4e[�xV�J	2�܄�`�n� ���e�k�?�?sj��.].^k��tğ�v `A�?N=I*��k"��(�1k�SE��R�B�d��9�\d����@�8	�-��q4��	'<m_|c���Z��|�}�}3\�X������ D�i@��a�W'ǚ�od�����A��ALB31+�Is�(�uׂ���CX����� q�GD�bע!j��G�z�J�|gΞ#�T,���'���u6)�EQ!��VB�Y�ߋĪg�O�KQ:!�X15���(oY��FՓ h>�9���]zy�sSɴ�Y�37� `z	�X�)EX͛^ZLN�\Wt�lV��6�}�/:��c���I�w�����:2nL�èȸi��ʷ6A��%����i��e���Y��_���[�u,�'�M�Qr���V�)Wh0�nk�6���&�׋#ߘX�H��жY|��`hB*��j�RFp����d�Y�Ż�"���'����Hg,�7�-��N%yn�S "ol���{o�F�8b]���j=�N��Մ(���[!��|?p�F����Cl�b��@��NBX��B��=M�.A$@�'Y��ķ#O�(�8F��le��`k@�G�V�:?BR|��.�5>����Ӯ�`�;˲c�&?留8|���n�=�k;�Y�=���`Iаk}ۊ����9x)q���_���$��rP�TU�H�/��RO���~đ�z8	� aӁue�ܡA_�r&�g�J��ܣ����"1
LU<�Sۉ�5��˶��,j� ��8�<��{S����Z��Sκ,(!P��兮��b
�FV���Q#� �
,�W�8������v���(����_�������x����p���Z����"��[e�?,��}����_�9�FM� �2�>�T @�1��a�Ι�=�π���(��@��8��	#��A��P�p�|(�����sA��|��S�� .2��OV�s����P���
�>�P1W]����?Γ���l���U����cX�U�C���J%6L��3���a�f}W���;�&�`:��]�eYX��ri%i��>;m�8��vM�T�����2<�����<�暿���3c����M��H�<��@�&�}�\�ĭI8N�����D>�A��S��PA���I\���6m
s�gO;���z�h?>�KCJ^���\w�L=���\����Q�{��؟f�t�;� ��(���\��~k} �kM��ٸsQЖ������p7�*��9J�y��[������
P���Qf��Q>��ki��R��1�h�d���"Ku4�[�5����G ���Mc��ŋ1^�x�&7��,�DwNFF�y+_Hf�%Ƣ��[��q�j�����V-�Y��;�1'ry�?6�x�����&�Wҩ�"#�Ĝ���
�T�U�Ek��ï�'�������ul�_G������D�0ṕkD7]����_������3�Y#x���Ċ��d_������*���!�X�_���aZ<�8�Y����9&V�9�Kz����VW�O���z�kj��ϿԂ���m$�޺?D,����f�{�uۜh�P�}ݼ�╨N��>�RWjK�n^i�w�YW�H�'�	�\��i��"4���`����N&�e*A��B� 2'%�L���:��_�����s����1)�+�_~�nl5��|D�7�^�E��p�4]W�`EGm���eԑ�{�f��Wt�f?!{��>ߗPi��h��q��fX��v��v��j��e�)�w@��S�O~p��m�b$�+�i�>��%. �@�2Ղ�=���A���v�vK�"��&��Z���$�2�:ؘ�*ĬK-��Q��[7�#N���>���Q.4��q��]��ޢ�!�����Kf�l��p�o��0�,�� �E��v��/��}%�Vޏ�ȃ[Q��_��PUb?�s�g�\���e��.$�?BX�1?�m�|]"�3!�R0�TR��K�iBC�eHX_f_j!�!�J�l`��8���L����Gs���qc�oxQ֬�N��\�y���Nx�j�`��r+p�fj�t��H��$�zPGA�T�8��;���Z�B���}㤬3	K�n�#�ݮ�X�l�MC&��������H	�����}�+q/�Hx���-q���Ce<+�X��2�����n�&Ѣ6G��2�5�ח7k�9��C�ͩ����ɐ��/����*��Yh�۽�o4Kh�"1B���7�LGp?���z?o6���ح�И���q���F�dxm���`3��q�Z�R�:����"����~{Du�[#�P�#2?{�_�*��AnѶMxS�H"�Z�B��C�&�?��S�b5�D���>���WQW�[uLXiC�������<Ն-O	$��/F�՟P|�kA��e
Ҹ�M��]����x橆b�T��C���021:���-�����Ao2jc�
�`bR~`X��+N�N���H|*�@�o�ݜw�:2:�vlV��d��l�k�@=!f�G26I�QX�/Jra�����{6�4QF���^�����G>W"G0zs�qn|�t�C"�/"�1ˁ�`6y��6�����.,��[#�Z��D�����>��5UQ�ذ��-e���l[+S^�|���A\bLπ�P����S�O�5��Rrz�_6's?���jAp~�é���cC��7Y�mCU
�Gd|٬�/~O��ي�D��aˋ����CH����J=������W5�E�f8����n�ѱ������)���ֲ�w��*�A��'qQ�w�����R�x�h��#?�~�7n�����ٺn
4=&(�̓T��O�!NnRh�ciƀ��X��ÃKP�h��Ԃ�Ǆ��"�<A-�DФ���g1���%b�1D��i�����b�[���)~ݸ��	 ��o���R%��اv��?��s�����]dJ���g0�y�/�>�R�&'���c]�+���fx��j�����2�pq��q��%贪}Ra��H�ӿ���S/��[#j1'N���`Ǿ�:<L{8

�>$�����fzW�p�:x����8��\"�Xbo�%E�/�qz)�-[�Gp����6����FeR�ì����Z����'�YK\1��n
�����͜"|���p�p�=˫��~�Xz}Q&�	�m�dx��hL}zq��3{��빞:fPy��h�U��y�ӛ�i��W�!�b<�.{J�Uٜo'��(ة@��)�(�i�i)Χ�z)�zb�3�5��D=1����n��>�/��j�����f����M"Rg����	��Fi���d� � ��L�����SM%�61a���e��]�%=�ɱU����?!��Z_N.P6~=�u��^�o�X�U��%����M�k~�/K��@����r�S�+�����g�v.�z?bQ���q��u�f���b��a�����ݽ��xi�n��Z4�Rmw��.���X��o�ˢ�kM~�_�9+����o;%i�f�Gx���x����*��酢��	b�v�s��k�[���9uگ�v�[���&"��}>�+�?��bV�cE��ψ8��ao�D�szl�V�T�:�k��o-%Ġ�1I��rc�����آ��bKaM�Ye�R\�kM��u9��1+6������p����~ar�b��U3�=�~�䓬�esΝ��{{w����T�Ǧϰ�}EJ�b���'�[Q�σ[ҵ��M�4�l��߶9��	֪6�p�x/.3g� ���_2k߸��o�k;A��P�C;+����KOn���'/���mcN�T���4��t���!'L�L��6�R>�E*w��s%�|�7��[v���{J��_{�XX,����f6]��G��o���Y�m��5i�D��LG�i�&6	`X�	�B.����]��y���)�xz��ܶ־���rͬ�7w�M�'f|�Bz&ȹ�(F��¾�)6������E�ej�J�����g�������;b}a B��:��\���?�ɼK�&XoBj�g���C��]P���H�G����ǁK6U$�\�
	/�����3���a|m��B�Z�]��:����c&&�X�+��NOd澇.t?�u�R�<����j)PH�Tϲ�$��a��t��<��� ˿�d�� $ZM J(*[�
�9H�Ge���@J�M�Fm�X}k��=x��k�����F�'�cg
�1yR
�����"W6qg�� ��a��.�T1s2x�����A;�'��h�C��ɬԴm�*�B� �2C;��ѶL]�Ƿ�!����X��C����d->~G1�F���/�@�����}�Ot�����dj�1:��@�4�X���Չ��{bJR�D=�	��Ʊs�C�+��׵d~���<u@\ө�q:��s�xn�0���^g bs��}�d)�,X�t}����o0�����k1�W��k�[�6��0�V|^����7��2�����l�_�F�]�/0B<Zǜ�S�/ �!��5�`q����o#m��c���-^�j�r��-3<� �����U��88��r����ڱ�m�n���ffOA{�Ԅ���p�>������@p�S�X�T�&�*	�vZ�&&ވ�3y�4<���[f�eW��������&����^����X����d��;ʰ�� ;ݠ���� ��c�����;���rL_�G����6& p��:S�d�_��<��e�MH�~<f6~Q`����f'�ʳ��Cý
����4e��aT�v��*i�p���NB��ޠ��@N����h)�!s5�:�1���*o��i�%���uS��W`ʨՊ������j�G ��sF�I����we�$��d�!�Z4�G �=��HB�+\<�진f�Ob�����y�@\pMr��0ˢ*�#A\�#�^�3�D<�pkY�b����PW|l�=� @e)�~���qG�;��m�'��p��_��ݧ�����gfwd�Ε")��yj/z�l�k�,ܕhň���=�5���C�2m_K"f�ըR�f\��<�C�Lb:u����I�q�������������@'O�/{+�᮸S�Z��F��u
�b���g��� ��r�Yq�[Mr�J�{^��7�h���]���C̬��V+'�ׇ���I�����m=����n|�#*���C�x���"�ȆU�����
O�v%����4�����M����f��t`*v,"B�Z��NF�̮Q+���i
��fH��rǫo�p1E�[���k�$ΫoY���Q��o���Dh94kR�s�~���K ��G��x�t����J�(}G	�?v
r�^�d�/�lа��`+�$��Q�U��xm�y	$,�H| �yz;@;p����^xI��a�_��^s�_�D�{X��^�1+�[��0PO�>�ep0�;�S�I�e�o���^vj\�RŬno��_p+=��aT�7i���ҩPt8�9h���`�FW�R��,0�9���wn �é�����-Ŏ��P�1�v�[����C��)^����:z�'�_�dH�V��l����^�K*��S�z`�ṙ��8�PQ��	�A`��3{<�(����������v���l��>U�����>L>�sG�.�{�4�V�z��V�;M�
|�§͸��r��K�/��o���M�ד�U��N�����po�_�����4���.���?mR�-^�fױ(����Bk��u>��D,���?�
bY]��F,z�Q⢎��B��D�F���q1�ΣM��+�\h���B����"�ܣ��X�q���oL�.Iܨŗ��ŻS|�7�!�(�g� ��)�I5�ڦ�O��H�X���Zq�u�qA�Q���0Z�
& ��q_j�J뗇�~�AI�a����IY'�"�5a����n�Ϥ������b��~��tCwȞ2�:��S��S��_i�i���@�Jߍ���Y!h��N�7������Y��
���$u+���@�w~W���AT��6S/c���l�"X�Y������R�^�������q�}��&����Uw!:~3���R��B�O*m�'�_�I�Y�Ib�_�T��F����X��@:���O�L�� T~�s�Sw�q1��b��YT��"ԃ��r*�s�)��n�5Cq+V�,����N@I?F<9�lҹ�����t����aJe�D]������|2Uo)sYO�A ��������� F�y�I�I��^"��Ľf���m1 ���q��S�%EUOZGZ��F�;�jkpωP�%`I�M<�	hjy����#ǉş�@m�}���쨊��/��>{�.�/&�7�Ԛ;o�$��� ��,E�T��k~� O`x��J}�f%�����;z�Ol(�j�t�2�|I�} �d4)4մ4�;Q�
I�3��9}'n:aXex]g�d�mNT�qx�����;/eV*�Y��� S���+�C:<�V���.@��Й����������8���W1a���q����_}~��`��>|�6��׎U���FGY�1O��h�VwT݇��ȅ^�b��o�d#Z���0�휳E+�� q� i�C��}���p7/<��]{�+3�F�ȼrG���s'������&��jAH{�߶�G�\2����0�3R|(�b��TsJ��5�Es�c��ir���r�:/�m�y�J�mS�jJ�|c���F�ޚ�xV���;)vE�f�8J�*o_��پ�s�1�)�[͍�DK8��<�*�H<y���W�c����<+�	��a��� 3J��S�(v;��)��I�rL�&�����U�)DT;�%C�%�7��j�����%��9����r�P�e��b+�j�����}x~�șH�&�AK�MP�u�N3tk��R3Y�Y��~��=3.��?c�$Un����������~c�A�qw����F�h*���.]�������z�;���|�P�P������I>]1ӣ���t]J�$K����ᓑ�%*��f�-k�f��H�0-�':Wlf��]+!��u4����ڻ>5�ae�����F�<�͜L��1�o�,��.;��S�~��3�<僦����@����Ly��w*�����Q)2"d�y>��4apG4:
��O���F�� )q�0�̄a,�,��ͦ<�?�A󉟑Dp������oĸ�gLA�>Ȥ�Fl�X���{{J���^��afe��]�	j��l��E��>E����h�ڠ"S��u!���s�*��*��LZ4S��O���݃F�pp�:R��B�E�{�*L|�lQ�}:S��0�{ǂ1����$ XF���ђ$��`�e,ś�Q-�b�bn���S�cFDʼ��ĐE�	��x��wX7`|�����~������Y���Y���i?'����K*O�澕~8᢮��h_�I�h��8>y����e�a��q�.���%ts䅚�VִTb.����v�e�(PbL���^+���[��s4j~N���)����Uś�����x�F�������o'�������[��|%��N4c!������p�0.��ɳT5� �Tb���Ý�'^�A	!Oq����S���鏓V�
܀s���V��D8�P��-�}�����\Չ|�O	P7�g^�_}�a����,��w�E���i��"ˋ����/*�����$���L鄅���#��nm��b�yIb���L��E�������Spmƻ.����5�$��Rb��iA��c������
�Qtw��ʇ���RP��@q�	K_����K�յ�b��H�S솖�̀���N�=:�0D?�.���(V廜����ʁ�a'�j=�1\�j�$�@�l�Q�ݙغ9�lh���l�U�V-�����9���w����/�3���ܰ�!�O	i��a�HE��_��u�#�-E=�����D+���e|�Fw���R�,� C)͡|�X�ǹ��V�zʂ�`����D�퓦:�+hӬ1�����?��E��K͌�W��R�@1�R� �{k��ܼ� �KS-�����Ȥĉ��uZ��1�1�E�
$-�]����ϥ��V�	��1�V��{�JU\��ˑSM��9?�lsw:���6�Z�%�W���	���q�Po=L��ݼw������\']Wq��/��@�%��\�3F�l���$��pHQD���m#��Z;L�n���}/o�}؋�8�ˡ!I��l0�DSuv�\Ϯ�Q(��/���*:��]?B��|���	x|�ꉋ�)���-�|噍�f	�����T�E=�Y���;���3|�v����õ:�R�]7)��y�k�F���1�@K3{%��'2+�0�����~鏏�=�,�&�qkm�Xy���*�r��w$Y�3�������J��]�zFX��?i����a8�X7}yg��ϐ�%L[Yͧ��ˠ@L(1�]R8�}����P8֋��<�7K�����B=	���{��!�ԾD	�ɼǖ����LB2J2���ƻ��:�'�6�;�@-�ncw��♩D� Ӑsʪ��R�:�bCT�Rӛl^��X?��O�U�7�+�x��Y�Î����=S���:�'L���� e��=D�T����s�XT�c2]�]������@V۲͸`�o�U�&�eOy_�D��J"�	4�YaB/�ހ����0el���x�#@���԰�ЃfZv�LS�}�p�	���@ؗ���"t��� �;3Pu{�F#���;��1>���X��@P>N�"��ў�8��&�3�Ej�^�q/��v�پ�gED3�3c%��� p���7Z���o:��	M�m�单��p6ٗ�m������Ð\F�F�-U<e�	�L�{������1����M��;�II� s@����W�g�f��@����'6����qǹ-^}������(q�	�j�P}���̥M�� a�����[ݰ�6�i�ڢ�ƍ~��|�H�޻?�m����.x�Cѵ!og��;]�,
�]���My��Pd���#��Xz��/F��
/�֕��B����^�bcK���&����M�5�4ԩ�*T	��ʼ5no�R^��Z�.��|R��%<^�`>��]U�����P�8�e0J�٦s%��{�t�\��f��J��8��d$*Yu�8��I�%�����6���=X�o
��{�
H���*���)~"&������+z��61�&S(��N�k�b2�k�����
=�*����\̓�v��>�X�y��WrK�f����{��Qq� >��{m�⸆�(�_��ɪ��M�$�aDi£��7<�IZ/��;��\������IAc���L����0ӹ}H�]������|~�Q�M���n�s�y5��N�U�HV��yW�Y�#ݼ��FZ�Q�a�bGd�un���,���I;�X�����0C�&��O���<-E��V�$��
�j�"D�Z�X{,i3��7MS2����C'L����"��Jj�q��8���)*���e�BQ���+s`�/�X2��S*�s����d5nO�-j�Ck��f��$�lE�I��� ��b���S�zE1 _�:�V�����n��#�S6�"
��5)仴Hu�5�~�9���������X��9�+}!vXr,�n�!��N��!��en�����S�l��~��\W+b�?_q��+ܮB9z�X�k���W��I6�v����{��g��Չ���r6�wv���@aũ���8�>G��Ƴ�
��sGs�ѓɜ2�/��G_��E-�?]��4Q;©x	����1�7��80|�%ůg��tbk�?rp�\x={�3+.�Hf�b�4��Qv/{]&�MK�	��r cq(I�9�>��x�J�`!�+u�"�"&����
/�mKkZL42"e��e�,ģB����מ�v����Pߗr���+�~�е��I�w[g�����T3���L�	��<�o�����}gͳc&��R��Ϸw��Z-\���{	���Y�u26q\�^7bBg��E�O�V�)������p�΃����k{j��|�N*N/�+�%��ϓfח;��{m���D5p-�EB�L�j��.{��[�4�M�l܁meĀ}��"b����s�N_�/�_m����a*S�2K�q�/�����R��=�9$�l>9�P]K |-�+S��U4.�1�g�,��-df�]>&�%�{>�W��&Q}@1Y�"�p�S��S��/50P�q�j)�ٍq�w��p��ǚ�#��%�s½��.gҫ-�u�T2ř�窩�,h��ؗ�v�����d��+��}-B	��_-����d䌉��l����\�2�GD��_���Zo7LF�*U+��%3����@�Q~I�(�֤2,����[�����=�U�+k�֗��!Ƅ��"W���"��w�a���5����ӫ�>�b�x���E���>���@J�%���U��	S$��s����:^P']#�<e+�H(��3��Si��DE�Gdo%�����2"i�U3+���.b*��K�bˈ��x[�$�!��U�a�9�����O�V�A����@Zr�Y_���zY}�� pp*Qqm�5WdEO��j�H,�{���+�����u��&Vr��v��倭6j
����$=�,��P�s�7 <�Ѱ[ھStc������Ƀ2"J��9b9d�� 
��%�х�
S���۞Vآk�r�r�������0bt|ȗ?rZi#�_����!�7rW�LZ��ap0���#��=�h���qS&8�r���ۈ^��gOr�	=�g� ��٘�,mƚ�Ke����0g��b���V�4B'xl�-:�Ob%f>�C�+]ƅ��R�ˀ���~��i����v����.13��s��i
�����u�{�Օ��_F;F��4�5Ƚ�&YV�ѻ̕oґ��ں�ѯl�+���'�]�o8��`����f�M��$�٪q�o���C_k��-�o���u�W��R��\*߻�%��!����網�*�!w�]W�	��|(Q$�k��Ŋ��w���e��ŕ�	2đrAz�$.!8>�yN��q��>���]L�:�u^�������:Ԧj\A&�9ьɠu�
�-׮U�{�UG�*ꃶ�D�ĩ��Bެ9��<�2q7�qm�V~���m"�΅q竔	#���H�[z���'�?�
�~�����Vp���8��+�N����T� _v�4J7��qJ�"m�#�B�u�)Ĩ����]�>�^tL>H]I�m�Z�C��ί3��|H�@� ������LZiy4x�l���h�/`UV���.��>�%�ƗY��2�oܬN�o�(\������p���8׽.'�b85S7		�0�L(Fq;&�Ti���C�X��Lj�\�G|��
@�������$��&��������!W��W�q���CD������!���S؄�� �!oM�0��_�qBԑ*�0��+��q��7w���+I0Y���.#��|�KW>O(4���*��l��$`F
?~YP����X���4�t|�@Y&��h���3g��������[d]�ۄ��-�wsZ!�9����<�鬚�,�$�ۭ���8�O��l4ix%f�E�ۢ\0��p�p���
�H�ĺ��n6��D�W7E!�PBJ�����{Teg���K*_=��?t���5�<g_�L&r=m���=���r�On����͗S) iPW%3�#!���/� �z8�}��T�Hu
-��4<��?���o�$�O��U�2j:�)�Y���f�>��*p�)y�HPݮ���oF�|�n���es`�8�ʡw��sWy��a�؎�� �q�ƹ�`��
5D+F�Y6r�N7ui������ʛrxCx����u6u�`�Ii��z7�F?&s�7��Ӹ�n��`@;C��D+'/���K�'z�+5�����@�R�S!2+���v� "egD�ՀC�{No��^�y�	�Idf�hU^��z��S�H�8,1M�%ͯVbO^i�%C�O���2���|]Zo�r�ϱ��R^����M��3%�7p���JƎ�:P����mO����v`P���	���9F/=%�_n��~�䪡͊�1/-V�I����Z����gw��	���˔��P�s[y�S2zç�*�����X�j��9��ӌ�jI��(g^f��>�/�|1ė�{�����7����O����T�d=�=�w��ã+�]$lZ���2����2��g_�BȉE3���{wt!D����d��������.l�!^�s��u�9�b4z�kmZv� �w�- ��6>��;<�`�VDX�|ΌX��|AoJ}V��T�X��ۧ����)��C4��!�;�C���h��j=�44<LU$>�8�O�ܛkBC�|oy,�s_�G״������K��!��]�8,��	 ������]ߒ�y��W5S;Us�̱���9ݽL*F8u
R�c�.H.�h���Y`��=2"���W�,hh�������Z ��BM�-�q���ԡ��<�������ۋ�ݬ`R�o�`���7X�4ނ*�S�`��R;cQ�mB���H��h�{-y�y� 3����jB�]07�)60����%m/BхСTc�ԛ��6�:$�g�|[�Bn�R耠H���:��88�?��i�!�c�ޞ�B�?Z��Ю�A��6X�nˡ,��6�_����&q��󰊂���!��}yC�=F��.-i�#˩��|4G�����0��yRi�?t&妇��:x%O��q&t�i���u�I��i��*T�4��z.7K.�	����Va"�lj�Aɢ0���� bH�Z��h��f5~of~��8�@C���!�N�J�n��Ӻ�w�.~�v��5/���.:�Ա1�Z�+ڠ�?`S�� �v�Cݗ��E:��,�mt-m�R�y"K*���������l�'42����![���T��*�.&�Z����J����������w��b�?���m/m��q��@Y��+��n���'��e'��<��nW�K�Xc�CK��S��}B���.[>�q��gFk�W��#�!#1�ٚC��q�>�;ҽ�Y�ج�E�����2k.>=H��2
vb��*�>7�%��2�	��2@o��fG��7�//%�yGW
r�jW���~T��Jnxoxd0�A�(_�,���ݧ�j����z�ؾEA������h�][��w4 ��}�,��mM���no����ͺ�� ���ď���c�cK�L�w;�ʆ�A�՟���vSʄ8�Z��s��w�]��>.>;b��U��v��n`��-�zac/QJ�|�1��E>Ԗeu��%���=�."Jun=,U���[B��U繺�έ}\��_�l��n�d�u�(�8�5aپ^�ͤ�W8�e�Ü5�G����$'R��Ow��u>��ñ�z��ng��k�g��<�T���}HWpu�wJ$���:q��tBe�]v�9W� У�}-l���Gcُ ��H�������[���9�X亝�����u��V�Zy�
��	P�^�l��RB:�BuF�� ᕆ�H����~����ʞ��p�-Q��M��'H�)���d.�s~���?�R`���>���Q�@o��x�`E}P�.�iu�ab�+&3������݄z㢪��qX�F��!��Q��;��4�O��Tߙ�M���=r�O��)l���~� �.s/�?��ݓ��G���r��x�7��`�شc�_�M�i%�d˄i��:\2s�� $��sڎη����B�����<��I�����W�/����v��6����.1�:'N�1�Vڷ!�o�b��͆5���� a<E��S0[�&x~P5V��Q��غ�zO�zN�TE�qcVݯca���f�Zb�(�)�a��&�]���V1lVg)�W����V����aVcT�5U�ֺ��6�E�F�F���2E�HJ��IWx
3aT���ڞ�fvQS����3/����u<kH�x,��e׮�x�T$��Fu�j��Q�lȘoW��R�%�s��`�VyH�>%M���I�WD`ty��]E k*G��%q׼e��T���Shw����av�8�>h۽R=��^��H�~�2�B�b��a˽�?ˍ?k����@�O��\�m"�p�oz����=)4(L}���[�5�gmm�h�Ehr���l��> �M�s�����h���d��!����I�P���f�B4)g_s�����H7!��E]�b�O8<?3xM��]_<3���	#����h�,Nk6]5'0�MzU�����/'����},�˧��O�D1Vw��͵�G��8��)#�Ѳ; �5�� ���^�'����"��%�o~&��լ��yyEmA#e*�1��h����|�B�{`eM�J*Y/F���tis~*_
�J�~�l&���=��Q̂��
�[����Q�u�(cL�{'���$�wġ���n�.� �2�pZ	��Y�P�r����N����-�*�\��d�/q��om(��F��J��/�Nz�=�-YtT4��?L�`&Ҙ1Z�o�N�n��:dr�������2�)���5�&f�N�2�� �*e`c)���AY'����A��Nt�R-�_{	i����X6_��G����,`�3�[�c?��SF�}�Sà@���&���PF"g����޳�ͺc# V�ި.�?m���8�ڦFed8>'H�]�]^��D%ㄏ.��բ�rK�|�`�g��e��9r��ӑ��2��C.��XS���Bb)�f&����8L$4�$B��O��S������s$6��N+%k
m�+/����:Ӱ�*- Ã�x�q�pZ�4q*��;�M���ۭlTCL��D'�r�7�9<3�}O�C���ዖ�9O��:]�k	�Vj���m��� &'��wsW�"���Z��R�.����]����ިU7_S��l5��7Z�'ⓛ�!���}���C��?�Iz��?v �#l���beܐ��p���)hoO!�l��7л��E2c��w��=عe�
���=�C�`�s��dl��=�ҷ0Pt�^b��>�"f|u�69�Ÿ}�(l���?��K������HN��;��[�׊�Q����yB}���ˍ/�;t+��4��|L6o%���,���S\��v�!��I���Ēb.ø!��*�O�ڹ�E5���-.[ٌ��ܼ���蜮?�]�>�5�(��EY��X�l%���x|6�X�c���|���T&�0M}@����7��6�R.���6u$UZ��d�7Ok!�w��2��5��E�##m�Z� ���FkK y�]O7���E�Ո�@�B��:�]tR�@]�6�"҃C���$����`-��yj�ɿm����~ݛ��������hi�a�2�T_�^��Y�������䯂t�顷AA5I[�mb����� ����� �	~��'z�X-̺�n���N-)ٚ/�A�s�������?��q6tp����($t�ǲ��&���eN!P�6�M���xO@�8�$qd�����`h�o
LڜϮD��3+�b�����w;�f���3���ċdݢ��R?��K>�&nG���b�*l��Yi���Zj�龾p8�����7��I|�����*��J)/�B�F_��{��2M��v}�H�@�
�iir�<��h�<��AT�K�x�-g:z���Rtx"�5��
~>�vnco_�5&����xDs/��$h���F\�΅y������5!�6X6�>5�(
�/����u��҉	E���~�rB>"!���E9����G+L�f�KDII�Ҝ�g��q�o0��*?u=翆�H��[��V?�I��s��u���?Rq��&�J)��H���T�-�8.eo]t7���9|sbb�L)�����'�N|�e�M����؎����K��D�a��<m�L|�)瘈!�+_U=�@�QѴ�"P��q�;u-{�_�u���m��h�[��eR������U��a��L�u�p�/3I��3le��RFZ��rR�4q7�c?���w�8T�˵L�~�@�������5l>�&]��|U�-k�ou�On]%Dm�c#�^�u�>�4��i�p�����Z�#�]���$_`h�J�ց�_�q|a���������p�<�<H��eC]��xdW.�3G9�èŌK��8eO��>i%�+��q��Ѳ*��8��9��%���`���{Qݙ��f\�T����1^���>m��h=�J����b�y ��s3�į���>���αw�q�d�)��-|�A�d�e=s���SZb������Mt_�H� 1j�{�����յ�Н�Я`qMD�}+����d�d�^1�@����������|�q�u����V�S䨼�;��&�,��?~4Q��_g�q@y&zb�L�Y�<���g���#GuE��������i�	�*S�����٨)(�wz��'nB'w]�n��$��5��	�0��‍0��O�����1s�?-P�>�.E��E�XqNL�=�'/㍵�qW�qt���Q����a�������$�3�4�ټu)����b%l�K�+V޾�&�g�6n]ַ�ӳ�1��U�����qE���?���������@��(����u����2�'cvZ9�/�R7���*�f���"JI�����#>];�/�>�o���^q�)D�J����mO��/K?�^�i��4"���d����u�Ҡ���--�NE����[Y�,��{a5��V?�p��]�eV�������M=�o�L0����+~�O�z�5Y���\��"�������ֶ���3_�g��qi<���gC�v�s�$�qM���3�T���R)��J&��w	�G�`�7����R<��N��ݤ#;ɪ�&��j<lB���Ƚ�	H��y��|"�t�qh8NHA}#ϙ�Z/Q5�{6Y��Aިǫ7Y�l�H��:��d����K
I� s}+w�4#���"��c�*>>�G��}n��`���"��A��B:���PO�H��)��M0� cQm��X�v���5�N���Ȝ��H!k�2�vr�A��ϊ�?�\~�ow���W�pD:�}��p���u=ꍇ�h���TAA�$��P}oR�յ���^�,�����
`��������s�Ը����ټ��!M�}q�����[xAG�Z���s �V�/�˗�?{�}s�'fOSTm�%���jeJ���
p����	N,�����ʛSaХӉ�@D���(���SE�{�R�˹��7cb;�`.�_��Eڕ��B�����ҽV�{���Zw-��;��Ƶ�F�v�ݟ&|��֕��(T�J(�&,B�d2�H���eJ���6PR��1���^���H��Mt9R馀�G�WqұS����yr�Y�@�x�c�G�<�+� �P\T���7G����B��<qC��}�~ۍ-$����_;�\��Y��>�J!�B��h�ge��Tj��o����+ϒ���K���sOA�M��b�߇� �i��x�
�	����X��
3NA��XC�"�ˊl�z��W>�@����J�R�`��㟁��z��T<ҷ@��v�bM#�s�	^q�FA�ߘ?x����6���ո�͢�1<�d���|���'z�ۤ++�����~������� (�+�r�~�T:�X�tc�R��ݫ`M�]�ao�-ɵ�)�&jO�W`�֞�!0��v�(��kWCJ���M�����W��f�Y�uw�R�5��нs�^�Q�{�X^-y��1c$�?�ר�E�a!$0��q�Y���A=.�����G2*��5���ټr�D{|=h��v"�&��_g{��׏x��jF`��>c��8�ς�d�{���_oC���u�U���s�`!^Ǣ�b�������r�P�컑�߶�&cG綥hyT�m`\+�_����kj����Gb�䭭=RAj�h�?u���	������s�:Y��\J9�n�L��q2����Ao����_��}�����Z�)�iU���` a�����_�S��k�^ƪ�Jf>��6yN=��5l�@{w���Bli���3�q$Ė�	壡��k��x�����e~�~�Wji.r��`��f5V��O�� OO��Fw�~�P��'6T�5`C���x������~�*0va�౛bjL`) rXJ�T�ᬬ�=X��0Y��R��b��B�c�h8�35���w~H���<"���2,�����LQs��W/s����� Q��¼�"�y	Jh'�:�}F@���)�}ʫ���Z���-X5�vm	+��"k��eVO��w`�'M���栁����|�X{�o�t�0g*ѵ�����/ �M�V��@�T3ʱ"W�N/d`N}��)S�K�{��E����e
����Xg,P'e�#���u��K�$�,뫤�?�����D�Z���|�|D+�,K׻F�%�Q�.+C�8��	�#�+8݈�v�P2x��~t��"�đ,릣:E2���)H�1�"`#Ĺ�U�u!��}��=�,;B��H���?͘�Ș�x�D@޹��k��G�c�۸V_��d��`p>��sX�����eLK/�kˑ1;�Lۯn��:g^-�����ﱦ8��F�4���\ �����?w�D6�w_\�1�pk��K~��'��t_��\&X�n�:	�x�b5�b�~�Fx�V6a҉���������d�� ?�FvU��x+d���H�f���&�_g��/v
���TkX��[F�z��!iu�}�*f"���6��{~���ȓQƧ4���a|!�o�E]2U�+.����+W�|��/�٥�yi�1�>��ނ�$�?�ῄY�G� �Gb�����6G%\�ޔ�k�OX�[�m}��p{�+I�����"�^'$;xl��%a�h�#0�X�I|�/��]�G��A١��(Q���-eEBm8�-��|o����2@��|�.�ɠ������T,h�18#��\�9Az�x�N�4�Ě�[�;2����}b<x� /��^���i�M�>��2�ȶ����6�)�e���ɯΝ=N��%��{���Z���NT�d��6������@�z�E'Wo�ъ�A��3�y�a��	�E�Of�Ѐ��� �����Ȅ�ٸ�P��^Gb�$��Yj�W�ҷ؅j����k��U��د�g��3C��G�A(�~9�^��Z�6����I���o�)>[��3�gr4c�@��je[�;�©���?�ى���p��IR3z�-{���R}�ۻ��م���vfMg�z��ގyP�os޺��o����?i�F��|v� �E�@w=y���zR1�S��t�J�6�0=%]`�N�;a�0J�c�+�����=)�?őw�I�>���0����$���Y����r�-�i(��{^mla��я��o^n>����&�U�`��h��ݶl��*݇lj%�(f�����#B�ѡ�d 澿}���S���6k�r��=�v�L�	 <+�M���J�m�:��FO�u-�II�߿��voc��MY�O����cIN1�t��0���I�\@gό;��O����c
�����1�D�J�Z�
�H1���_[��W8w\)&|ϳV������}<���.LP����=�Czc�`L]ب���%U��r���~Z� ��qC�]	Ɏ�>8⻞�[�"���-���F��x���	B'���e�am>1r:���k#���?�'�q��o(��q��w��^O��$��~Π�Y�72�d� ��`�=��U��γ!�N�E�N�F9�����"p�޼�(�C������e�؂Di�l>�xi�A� �.w~�z�`bG��OD���r��{�`x]��{�4Q@�sJ���΂���Xq,T���1�FĬf�o$�Ԩ�>FI�o�n���Ƈ�.�τ]�����ƌ&��]�E�iu�c)�ij�N�oJ.*$�EK��ju��e|�ؒ{��'��~��������co�p7�A�XA���������Ĵ��s�G+�/mth��g�w
>���I��>��)��J��wbqb9�")1�K�R����2>`��H �l&�h�u�(��R�B�P�4��@/�Z���AS1۝�?LPU���*4�b��wQ��y{C.�oc�-��dH<[�rP��hF���F?��	X�9*��>�RP:f�e�z�T�Mn�����#ҥ������T��f��}���oAt��qף�@bb_��$Օ�	Ĳz�u�&`ėח��7�D6��!�����W���oo����_=�ll]�F��m��ӆx8��^�����v�UQ�� ���I�_���	��U,���K)¿��m��2��5��y��@ܽZ��F�:"��s
%n�NQ]���\��2�X� X����ý��n�K��f4щƿ�f��U�����Ņ�iLN3��i����ڏl�r���	�h�[x^cH��JL��^�h�����t�d2�nJ!��TwK*t�7�����9Z!�P(�Zǲ˦A���3�W��s�i
w��5�N�ǟg�� c�Q5ǂj���KmgΓ�_~��9�����#m�[�%� ���G`b�u�����/XҜsޮ��b��+�xB&��B��J��C�2kٲG/G�&���q�4�`q^\d80�wA� 7�0Wۉm��N�g��oA&v��?[a=~:���Y���L?hY�T�V�'Ö�T��W�"�۲J�@J�IRd-��u�Z������$�PIT(����HV,A �ܩ�Q)�2�!�J#��Tڟ`��Quxh �(��LO�s)݋�?�OA>��۴�K��0��b�T�Ϲ"hM�(�q����O��pXC��A@�3�y�/���_�{���S��I�ZA�O
����"@z@��SS;��&G���'�U��*z"y�_V�X��ڌ+��T���k%9ϓ)8(4��S	��5&�� �N2��?��?0�8K��g}��,��HM�M���P<�쮵�zG����vG������64�!�.ۓyr�r���Z�W�P��?����7�Q`�/p����%��S��+���+�?��$��#|�򯰜$��������t��V�i�е�$_=X�^���S�D�L��H׎K��Տ����;b;���^� ��>�_��~z���!2�̝���G/�y��:|� �Gw[��<�M��h�4��Y����,c_���YȮ+�ꌢ����L�l 믬'�����Nr
�֍��k4?/���P�dhw?uj}Y��M��"�_�r?Ee.N��L�=?T�^��v�r#��8��=�=~$�a��S61�et�$O��_r���y]�ڀy��o����ﰩS�/|��Ĩ��Z]v���}-=�a�t
�5ձ���ԵxY�vl��.�_�����[4�V0f��v�8��֟����/'#�~L���Tf�G�{�ec�!P8�Q�����Y���B��O��,pE�����"�N壊6��65�$6{�~�2�l���c>�4^��(¢�_��+����ާ!\�d(�u�Yʃ��Ť�r%&P���� �zȰ?��َ\�uϴ﷝�� EsJlQ˷���/o��5'����P��6=��2ZrT��>�8Y��x� Ɠ_��e&�'�/2����,d����̝d`5����a��n)�ї��-��،g��P���k.+(P���?5qn�~�dc�N�].Gc�c����T�L�������%�\��
�T6m����arC9��\:P��.z{��s�tp �����	
u�ϵ����d8�� ?�K��b����9�w�]
�
�8��'7�a��C(L��8��,�u����f �T�9m�]?;d�F�&�4'��cf�_$)N��-��d���l#jat~�j.�JןM\�~�����/��1�� ��b3�8�T$a|)s��:쇅�DD�Xb���?���L4sAh�*?�����>Pm&\�����ϐf:VM�G��22T��rը@�M A*պҝԕ�6;�'��+��T Z2���-Ѓ_�Z���������K�M+�Q����C!Z�؝���Č�Y?�����h�Uk:����S�`T��G��yl�4^�X�?޻v��7�F���i�����${�K�,�m��,�#t�����s% ���W���C�O���HJ��B���q�����$�~�,g�,a8���-P'��F���Fd�W"��4+�r��/��%���� ����BWh
w#�BJ ���􂣭�͟��:��.�X�#��>-���?�=w���)\�͒x~tڂ1�'&�䖠2��U]bհ���c�+�M�q� N`�:WVRϪ��w����8N��2nd`R�E�,Y;�e^�&%F	5{��'S�J(���S~E�-K�c3w��I�g]*`���"�o֧��kO���5:�$#����	�a�"׏"����ͦ�O�� �Y4(�oPi,�W��.A������-S�k���g,)G 1_x��~3���� `���7��a5�����F��,�	�ˤn-�j�TO�
_�S=�G��$��N�F�A{�h�<��<��<q��F����\(o���ܸ�d��&W��uE���?V(T4 �vJ�=�?�=���@�&���|9��5J8*-2#m4���e���9��r�6���C`@g�OG-t'K��l��E����]0� ��4M�c�W���y�J08�2s#<�3|@���8�>�vF[�0׽[uh�NX�p��_�I�d�U@���W8��x���d�#��Y�S�p��-NQkh|)�U�MJ�J�RR��k `��"�^����㲲8B����JB���BL��m�X��o�B�!�ϑz����1�!M������͗%���Xur���-�:��J��|�]�u�T��b8}��}Z�7��߲��Ĵya��T��_�̘8��ӎLÅ�!�S��*�?���}ǳV�Q���~�P��K:W�b���o������j�ځ[Mq��-ݝ��8��S���+�U{g�Qr��v���r�N��zsw�[��yid�\�.�X��S�L;��'˘LQY���{r� ������,�LJ�	x3�0]R%iX ږ��Y]�%λ�8{̍��)�E��*�����Ч���+�K�m
DZ�-D��䬅w���|ӎ��8�b�0.�,�~1Ȥ.%e�A]��e���
��%�Ai7�g$XU��s+��~�( 9Ѹ�嵔;��� �Jm��j��J�MH��*ч��%^s�F	��8
���Gen�܍�l#I-JHy�Ⱦo'�J�'<���h�����rNj,-��{��A�do��L=��bT�?�Y��FO0��������~͐�<a9����6��oTPǚ�%�V�h0	p�� �
�1ʉ��ƶ�x"o`C�|��Zs�'6W���D~�ެo�NfD��X���_�0�w�ظ��V���{U8i
�ٗ��idn��xG�2{_��,��A�:c�Rx"wo5S�E��k&��.]�����f:,WG���4�A����)�꽣и,ݐ� ���G���(u������������F�����I�!E��{3=T�>���X�9K�b-w��Z��b?L�)�׀�KI��>Hkph�7��DSl��u1��nv�z�����$�;E8��f0㚌	၈VB��z�0	0^�RZ�_>B&���5y8M���Àl���&$F �� ��}1�Dx�&�Y�P~��P�L�#Q�������;�}�4��>�;�~���&Mwe�ܐ�ˏ52��U�D�@�;�u�'F_U��Xq샗Bt�3X;�Yݖ`:� 0��~��	��0�q`�V�����BŚ�3�+�F��H*L[_Pu�}?79�~��lo�xL+�q}�L�P7��A���\����sl���T��jv�����V��C��{���|O��*�y|f�V�������\6�z��j�1q�V����K��x�˚� �frQ��.7|�éoP��Nv�^��o:/	Rp'��w���".�DV��J�5r����/,��(ܢ'� �ۍ�ּ�0�Y�߄y��#uR`#g���G�~W����p�e��Â����J�GM/��A�P��^�l%Y@����i3/L��ݼ7�R����z����<R,}]3��K1xF1\I��Be�~�+͔��j@=+�Ϳ:���g��-��c>�t��~]U]�؄��9���/���vt�_��M���i.D͊d����T��7ܖ����<����
W�����s��As2Y ��vOQ=��m�>�)u�����u���+�mw�:0��sR�����n���V.�A��r&P����4�8Ws��o��3s�Q5�n�@X�:J�ac^������~�@� �j��`Y��'���__4ʠ6�[]���z-%wD��1XI����|}�HҬ �,�=\|Ǽ|����J-���,	��B�����_�@U���3�'"�$�,F�`�)7��1Q����$�����������}�"β�E�V�@�u��-Yф��q�mk $5$�1�H2���}Ԥ�I�$x�pq�2Bt/J�^�j\����S Xj�M��g$�G
U4@�S� �>��%�������g����� ���T[�lD�j��Su��~���P���Pq����9=�uIFqj"��mk��T׌;�1��	ٞ:�f��Z ;����B�a/V#���yZИ�=��\3���3�5�J�)H��^Y)��wLg~�T���(>||G�hʼ!l�H�d��1<����G�����~���X\1h��	�FV��CiF���dD�ђ�D7��(�H�����X����E��CY�ċ�QMi�0��:���	C�|.��ap��vj��t~���Ph�l"�.k�E|��4�k����_�`�� մ�wd�Eg�#r�e���d��<��dֵ�����ǲ@�jP������x���^�QF4��*��k"��~Mh֏j,˴e����
�-��?u.c .r$�Y���_IL3l2��r?����-��
�u`c8¤,� trW�\6�²�]R�\hf4;�"�.�1�����*����s���ІM���\�@��{N?��	�n�~����������������}(M��rj�h���[US[U�H��I�b�(h�mM�WN�	��ɜPC��94}g"}�Q��#v�ߟ�
�����8ߍh�}E1@��(��J�'
W��t(����v��R��<^ûG*���2�n��{�6�g&Nr���A
�D<��?��^xBp#� �Ҝ�a`�����2DTl������������j5��xq�ؼ�̷-�|d#�'�W���pw7�Q��j]8��y�HxR����o��վ�,���QUSN�0l3Q��']�ٴ�S��O����^5�W���t:7�fĨw<i��<4I�d��S�������"�bp)X�S
9a-m�C:�l��r@|�F��㫑�c���i:ib~r���n����3Y��&�Cʓ�-��7P�x�2o��31�U����\-��m`���'���	�:��#u�
��q	ń����$T�ЇN�~7b+���������V�f��CD����(��Nk;�U�KQº �����4�9�&�M��M#���_�i�����Y��qƳ�`*�w~ ��`�aBU
��=Mqk�A��`E���oM�J��GKO�fFj�&wb+Պ	Y
T&�Ƈ�=�D��[)�	7ad/��R�7�����i�m3����쳽P��R#���tC�@v��w�	�^�TX�V�H6�OV>G���͋�@7�5�U��EZOխ{��Y�Hek���0:{�p��&�_^ �鐸���>��$&KjG|X-��@�>h�[�����M x\0S���1X���vV��� �V'�����6�![�h$ ������V��r�/���~`�G�p{{^2��Y�:!Kr}��	��5�7J�e1�q��>����`��|좡8��jp�QQ^^���#��?� �����_��;�ԙ?��.T�2����B�$����\�}������q��FT<w�ɎU>f���%�f�)m�i9��vk3��eti�FE0šLbY��o��*#,�t�`K�����w�E�(�0>����9}W\����� ��P�"C��c\f�'Q�v�������BBWC:�6�>�{��͠�Þ�Wj1�G�q�鮓ݯC+�im� �Q �ZD��:���u~��عA_��$���myg]`l꧑`	F��VAz�����5���M1��9r�F�貃��.Ã9YB�IT
�]�:�?Yk��):=x�[�$k�@�-������0�z�e$U��mz�uFOZ.����L��цH�c�ľ�!����DxB�2��[1��`��>'�[�h�Ǚ�ȗ`���3�~��Z��W��6������̘��H�H����:�8-M�j/H���]��;n3�!�q?�>�Z͋���������MP/P�p�񬿧J8���G��X�q�����@�Ӌ���g{�Ȁ�.4}�X�5'#�{'�c�F����t=Ʈ�Vŕ��9�<h�?���IZ4S�ƀ�]�g��m9�&���9d|��R�+�Q�������WG1�41s�[o���j�*z��WD��
Ǹ!�	�<�������Г10@��Ƣ ��8��Zl���X�O#�V2����ψ�)f�h�2X����q,��ѱ���B����hWR�i�9��]������3��ױ$9(Չ)Zl�E���p���p���0a��&��S��o��!&���H��#=�6d�ypc-;F�W����I�I|+E�K��I�m-J|0|rW8��7'*S�>i�J9?��/o��B5�U�z����1��+tq��|M�T}{��b�"�*|^8�:���c�����O�JE�U܀�0�t}.�K�#�,��Ä��v�z���e�-^'z[��b+���N3�X��l�>;�EKK�GV�'�|Vq����(��َW��:�P��v$��,ҫ��mz�|�:U�4ZY6d��̫�d��G���2F&x폧����"��{������=l���vVoWO�Di�ÿU.�g�/�Jaȴ9s�4�!� ��y���A�zYy�0RRl��X�p9�|_h�J��E�&�ǧ��eRu��EK�TT�t<�=��(:j�Dq'N�#`�< ����4�n�j�R��E'Y��^�
:�y��{�����$&'p�+��O��X:���H�a�\3�;x�w�,|1��\��Hr��qA��������v��*��e�$j4ï���}���b�>����^n�"�����F�<t=����шQ��������.���=]���`��=�PP��W��(Ğ�]r���en��Q l���̵�����3G����w��Rq9�K�����}�UAxg?���a?�U!��k��<�A�S�?*� /-�:k�G�� 8&"&K���۾�˞;���"�/;��m�!��?tT2��y���*��`I��߅6@C�v��X�ڭ]�Ş�|�,��L�Ҿ����m]'ŝ�B�ͧ)����5~�|��{�1�{��!���u��ʽ�jr�U[�����l�,rE�v���r��gѨ���	�vkcW���~T�fz�hN-�m�7�Q)*0q�w'�`Q(���\3@�J�-[�僽lNM��4b�ߍ�#W��vf �1��q����G��uO\V ��5u�����6v�ǰ�W��l���W�t@��24m���-cS+qh��kܾ��ŋ�����	L�^�~B�.�b �5)�帑�>�>,���MK��C��|#��,V�A@%~Q/�3�׃A�\A-Y�?Z��R�,f�{��@��0>Y*�w�CŅ���1�T���U��������F0Ta��q��ʍ�o�����	�9R<���6��?��܄Gh4���0p+��������o?Y�A�T!�\�S�z�;ÕW*<�1l�����������Y��GS���~�<o�Q�0�R�f`/I~#����_�A�9�S=ROޯ��}s'ǱZ�ة��9Q�=�]i����O�E~��QK�i�W�-]��D�9Q���Ev��K .C�J����Z5�
C�%��x�(�����@����+g������ֿ�C�bB�z�+�a͟��18Ioa�a�{b�OJ��/_��)�p��x���q_���)�D���H�*�Fģ(��n��:��=H���u� �;�T����Mk�^&n��������	]���ع)�e���[�_;G��1W� +5�Q3}ڗ�r����XK��c�?DT���i���7nUoi�I�R�2���q�%	J�J�|��Tߐ�C�it�>V��dB�8�έ��y������S�L �.o2&^�(OG�v�(��eM��~�87ݿ�������5�i��2��n�g͑ ���;�ҁP��e��R��x����`�P�0�6Lt�-�Lt$�M���*,���ݦ�.�f9��\cƥ�{}]�ߜ�w:�u���Uڙ�R�8YY��M��v&:n�]���M�&��4��?p�Q��D�?��x�>�#}}Xo�mAN�1�#X��/j2�F�,�ʃO\��t��TJUe�u	���q���Pj��UOG�%�&�#?�*�]J�cWM/;e��.@�Á�gM����Y�N`95��	Wy�ܔ�:��	Y��&u�1y߃{J�'�2�O;4c��U�Ų�)p��B��驅���#��-�E��L3�M�{nñxQzz��˕��_����[`R`�� &U=1��S{�R�fc�9b_Ioo3�H�\�־��u�o��8��Jk&�;��L�-{R���<�[%;���?��9<���zc�q6j��6��m�vۘ��ƶm�jؠy7�������d��[�>g��Y��D���&R^��W� �B?R+l�Ð�w�u�a��Uֆ�X��f1���j�T� l�l���	��ʉ��4i��c�E��l+�)@�]V��r�.�.��3������:ibDtm*2ڷW�:�}��Q���lQe��Wy���˽��x�ώ���_4Q�(n�3���:���]�	W�|m_8v����"�I�>�;N�e� �V=��O}�=3X!���F�P�@MO;�@?�l���:�5y�Q%�ڏW���Oi�S�ZO��ɦ��R�ߨB y���j_+8�*�juLrj�5[�zԆ�퉵S0mޤ�Tj�C�vQ�\��������;�FŌlv��W��+%��t��_�������������W4�t8�-�L��P�!� X@�r {�2ב���v������yĘ����o���!]Z��~vD���F,��FN÷�$|��-�>$RZ�~��H�w�4fb��OD6'�Z�Zj?��@`�jk|��������8��f�{zNd�2�������E��{�ȁ_���Zč����~ =��/;uz��1�Ķ�9=V�I9���29Q�)7�J���7��2������ܨ�/��,�'�-��$k5 )4���?[h�=sk�yK��S��B?-��+R��wi��%��;��x���.��\�7,��Z*'ޟ�*o��,�1�2x� �W�4�:Hws_K�$��;����L��	��yK��v�S���չ���I��HZ�(�i��Ռ���W¾�_h/�#x���D��T�}�ǽs����苼~�>j���P�)���A�v��r���y�Jj�&5v<�0[ۍ����p�_����W�-m��9t���5>ˣ�"��X�;B������wE��w}ǽ�mŶv�8�4���f�6h�-��T����Z'�qJ7�,�s%3�S-@�wP��~~]�^�&e}�2<8X�;��	{AP	����/��=����Z�j�f����Oz�M���~s$@�~KA�Eψ�ɯ��`7��7�Y ��N�j����� 3���T����ᖻ�"|�x�DR�
�hr>��tG�DI�8d���	!u���+��Ȱ�8�U½)8A,}�W�Y����;h��5���aP�� ������+pYS���c��
���Mg]?��o<�����-�3���������T�V��k�+e��Ӎ�J���_�������ޔ�@)6�'ً����j��� 	�ɫ ����CN	��+�R$�.��7�{��������}F�׺����7�����u�����C�fZ��3*��Ʒ��*wO�Dw��v��
��� �8���i���J���]�{~ m��y�,���� �`2�O3`c�
�vsO���&�b^�=VmG��'��QǹߢQnS[Z��,��!M	��n;i��C�k��i_m�myG� J%K���w;��K7X��3я"���Z|�_(�x�M����3����uZ�v]�%��@�J�T"����,�!�,+����K���u/-*���t*��a%ޟ�J�[�v*r�G:/]bk��i���O�6zLiM�V�����t�4�mG!���Ԕ������_3-T'==;�Ϡ��%"��R��Ǹ��V�P��!��>�u�FS��bi�������}�k�y����u�z��yv�y�F��+j5tn[�2��Ea�n�,������3<N:Z�O8�\��z��_��KL��9/C8�/OCt�|H���t�)0k�e��r
\��_��?Ԗ؟���*�,�A�nz���y��� £�ص8��{Z\�����-�(���ӿ����d�Z���7����j��f,^`ÇL�u�2g!"����n��� v�^g�)cN�R3�V��C�/G��>!�A��A�z��+��1���ȿ��,a��CEC�^po����3�~��c�+�[�.�������͐H�u�ߘ~��X�#�
��Q�� ꭭����%D廧�r�7mSg����J�����A�t4���˂����^��Q�J����ӓ����;���fBٛ~��I֛��"�E=6X��~������m���;�Nk:�bt�[!{눛�T�R�����`9�h���,B�̻��|ғ]��;�/+���=R�cI�x�o� ����a+f%t@�;U���/�S�WTo�L����(����ٹ���N���[9˯�}������R!�?ɩ7�����-��{/�z\�/K�|��X��}	��eT���{搑�P������E�9u��]w�r7,C�Eqn�PLj���Gh�����x���Q��BxUVZ?�3���_\�ϭ!rT��'!���ż�������rY��у+��7��iyx�T3#�ӗ�o	��󰍜،�H��J�p2�W�/���P�x���ޏ(/M ��O��R���z9�� u�~���u�>������AK-p)n��-����t����6��sj������.:���*<�r�B���@V3�����4<���㺪����ʒ��m�H����O�	��u�� j?�J�|Y����`�l{{,��	<�U�!�&���RWKI�;���<�6����x�ʹ̎�ڂRK~f���;��s�a-d�y|3ל1�S���{�^�z0WΔm|\h�г��p���!��Wpat�P�ӭ�����~�][$������Hf�]�θ�M�-�}�Cw�J��e�;Uk��j�e(�
#�����Fm̧@c����=|�5ՙ�X��n�^���Zs:�W������jk3��ݷNp���~�f�<��5%X����a3�6�-�O������_��������I�f'-�a�r�j��a�B�x(Ե�5�~�'�Na��aG�6L<�M�N�O�{b�`VY���@�郟�V|���/�pѥ(�P6ђ����9������`R	T��/��स#��q�Z�B���9����ONp�^�O؈f����@�j�3{��HE-iL"!S�̫l�bס}�V6��3�ڮ��Sm:�VK�0�a.������<nI���M�Ӓ�f����sz.�����'U�y=�$-�� T:�.|0:qwbMN���Î�4��������y�g/X��������)����S> �@�.*p1�Z��C�%}�\I���Ѽ���;u{|e�U�ǶyÞ&u���)����F�m�IQ`�J1G� ����-�=?pK1���❮
K,)Ӂ�Vף	���������VR>�Z��n���mK�C:�g���}*ըz��9�@��̏Ef0��1_��1�j�.V���{�U�Ǫ{'�~V�nt��]���-� 5��ݒcm:s������~V�}3���f�؍�<y����Dy4�B9T|��Ҽ����69qOu:}�c*������G#P�9dRv�z�W�
jLY�$�6�RRR�?-_<�8���<��Ԍ��M)��o�K��l�N0�GtW��[`ќ�7�<*�"Bt�}�_��=��I;h�����Zlnd�@��	��r+*�د5���V_V7,a�>�^u0 ~Ճ�;^���e�]�q���������gϦW`��^�'�J!�Q��Q��UBV���&еD�r�P�����<'=~����cS�n�E�]h����C����B̊I^�P��[n��x�p\�b_�
��kcz|q���`O���X��e��E���E�iRw�U�}
7�5��Eu�é�n���0d�^�g�{G���-4�;!%̈́؞,2V�J���N&iPv�'�扥 �HD'��J�������){��W<��^��f�L����@�m?�1^�9:�~�����I6�;�\ai3o;//�k�,4�	���_֮��q�5���!66H�)�e��}۹�&N�^ڐ��_�u-���"�� #k����tß����,��醡�l�{O��}-�W�\��%�H���qk��À��Ο:���fB�ą����� �v�=3M軎/]/j�G��95r���t?%��{`�/c��&i����Ssc[,�(�k�%��؄�����MD 	���LL�9����q��]���������m3t�_.�[�j.�,B�X�Ł�����N�s��׼�y�)ׂ���E��Q�V�Թ_�=���&�r�fZb��Q:Z�� s��e;� �Ju���RPz�<��=r�ֆ���s�w?����-8�����Z�M�?e�����RdU��-�~ߣ�gs	(��t!��=g!�V��%SY�G3,=|�6X�>{��dSn�D��WNO��8�|g���qO�j��
UK
K\���V��G�q#�F_ �ߞЫ�4�
���{�*]�(�'�Rz�gqW���w��o��-�̉
�$�op��jp�%l�E*ްx�Er�\�=�J��"�����3��=B�F:�ʠ��粺��b��B'Zo��6�Q��{��.��%�	<mLZ��)w�@�_j~�P��W�l�Ѓ:Zq�+���.X�=�)��\�4O�ŋ�C�w/�4��,�y��j�7�M��.��>�x(y�e���o�	y�֛	GL:bt�s-����eM�Ġ�.�*p
�&g�	�h󳙶�{�ܠU�N�����7o��݇�����jOW�1��J�Kx/�����o�Ÿ"T$���Q`�C�`�̘���-j�%�`z��P�y�$�� t3��]ʜa����}�RT�E��2#C�Z���Z���˪s�ථN�:�(�~�,.s^or��o���_A$�z���+�S�N�����|�6Ƹ�� �]�zx/`�
�~����1iU5=�+����\��vbzS�_��a��f��ʠu%�8��ӏ~L��y[����9��z����I����)_��v�:������}�a��!�b��P�Gk�ބ$��ţ����%����
��f����b��w=NVa�2��Ȼ�9��v�ѵ ��ng%�r*��ղf��2k��/Dܷ̬���F��|&�ِa�B�n�}���\��8ƪ}����m3J�K�,�
T�<���Rv�K�e]&hS�_&Y��ś^r4+�{�B���?zХ���7ƅ�Z�B�P�n�f3/�1��b?>���P;h�2QY^�]�4rϱh��7�)�S3�v��<Bew���sm���S4�|�f�Vv	�^Z�ؽ�}�����5�~�_yݺ��la��)�D?�WD���9��l:��Mp����B�%���yA0ى��~�`��дV��A��a?9�C����8�I��҇섩��O�'ߺ\�|A�h	�g�ig�O'n��\��k��U�-�{O����Ll._ֈ$� �����n`�\c��^�`�_	��;K�Z�%�*4�B��+�FH��'�z9Ga7�T�e�J` �:9[��*�^��%<5�S��(���3k>$1{Rl$<˻�[�m���<�{�E��sdU쎱:�T�&5ڭ��c�s���9��;�p'��	�~O����#V�+���h��@qm��K�����8�̻�3�`B�{��%UG!�F�Ėee����^�~ס����N,�H����͒���/�,eLx�%�[蓼謚f��D�^�ƿ)�G��i�dϙ����E�y@��ʅ;XI�V�wj)�jc��ⷊ�����d����s�tuuݡ.my3�b�D��Nm�Z8�Y����}5+��x�;6q��q�|L���(�+Wg����+�/q��p��d�}�鐥�a��p��Q���WT�����*}~�i$f����)�J�8X�DҦ��mu�[�{1x5�$�y'6���{y��V������&�H��I��u[�=r+_����wfn�4��4�&��v��S��H|"��bf�l�b��9c���-��0�����÷T#�>�[�ʯv�6��亁�Hω�S1߽w���]}b����B��8�X&M�JG;2��5���c��������q��h�g�I����>6�j�fէ&\ �A>g%�O�R��>p�ǸV�HY�`����̶'̣��;��0p�#;׊�B���{;�X��f�E:�ٽ_v��ǩ�̃�M��_�yR̀1v��x>ܶ%�J�I �G��I��ۙR���N��.�"؏��h��ef��>Q���$�l.o�\`�3ٟE�|+K�nY@~ǚ��}��=;�����>�$�8H��.����~	'��ej���Xj>��~����x��{�\��;@�^�k���=�7��T����.�p��3M���N|�AR��LT\�54�
s�]�C��e���(+��%4�F���m��:|�(���Ѻ��;����n�����ϒ��4��|%�)������ϼ>�:.�h�㺲�ZͰs��3�j��������{��b��P�Зb�u�Ibo\F��(Ip���󺺄jv,*z"H᯽:�x�&��W���mB�EU�;����ݛ�"�SǦ�7K^��Cm��zw���Nx��Q��03lp��$��G[�1zn^VH�=���[F)�n�`q����qG�9������w_������c�n�v%��N4��Þ���w�3*9[�Gj�G�_���i����ι=�Q��5#��`ăe�}_q���� 7f�/�w<������k�r���>cC3�t�9���9�o��u���bϢ�1V]ahl�3�i3s9��N~�����){=�(⡮���#�~��*�a��F����M�G���Xt�Ø3�|�ǌzG�r�9X�͑��CN�܌�~�R	#�	R�xT�'@j�	������V��Չ���%�H���{ͥDB��8ߔ�1O���_~UZa�&��z���x�x
N��H��%���ܑ'���D(u{�b5�LV�a�����s��B٘E_�*]p.c�Ŗ�y��כr� %���]�<l�o]%�'��6`s����Z��#=��2A��>�e����L���B��@A5Ab?.Ϯ�2ĺ�b�P[�xs+'��R����MoIi�E�ͭ�C�/�'��@��		
��转��{z�P�o��,&l�;��W�s��0��-�3+II�A�L�H�����p+����"Y��]�����˙�q�T��h�.�>�{��F��������"�kk$�L[���$����>(�h4���gI�{ĝ�ȭrjh���ԡ�\
  �d%fbq�*���0VF}g�� q��J��n��I5X�o�&o�QC�A�0e����:����-pv�X4�uN�/l��� !�׃[�V��4G�R�g��r|��܅u���2�����Ȣc~�+`�牀P��_̉���WӞO��%���xe%ά{bV�X"F��&��%�wS�s��Ɔ����{�����pb��!��W�]'��}1�%Ѓ'�&aDBE�'��_�B�d�58�=��W|�M�G���0������x6���FHO����I�pUf�j�6�r��l,�Zq.���o	�X�y}��4��Xe5
i(A�A.f���$�Wbزm�[�J�ʤB��K��=��xȃ��w��;%!8]��qT������❯f��.�g}\��7�b��)w�4�^�}ї�>lh�
��R	V&�T �w�'gm&�4��Er�]�����ڻ��r�dh�f��D��a�y��uJ(<��z�Ո맶ȋM%#F�����xĨ܊��i����t��UB�� A����9�#���9���l	>��{h�����>��r�a���v���	g��� gg�{�/NS!oǇ�*��qY�$,݇,Hg!��U6)�kJD�na
%!W��C\wH>��ca�?��Nǂ���kz��� Ph9F��S^������c2�<y���(�-zm��q�6+O��Z�y{
]��G�j
�jD��'�ά�5~-�J'2�%2;�SQL��y*�.#��p��)qH��� ��bK�B޼g�\k�a@i .b�,�0�Nt�(�s��Dj� b(L��T�ʖ��y50����t��}#"��]�������1Vi?���4���D|rn�-��X�]FԊpE�x'ki3ڀ�fh�C�����(�W�埣��x۳�w�Ӄ:_��bC��sÁ����oRY��	)�4N�t��X-r�>ن���fP4[����E�Q����H}�7�&Xު�)��!�:k��,��KC�,�Hu	/����򀀌&� ��a�M��SY|m��y�ƮT����w�� �}J^�R�����Y����1�fΔI��K����M��œ}��d�.����ӫ��@,��Q֗�_C���b��w�a�o#siJ�i͂���S��'6h�ⱳ g7)���p�&/ ���`s
��<܎0w��c�p0h�h�5Qi_/̸�.N�v>��l��M�Y�1	�Q��u�/U�*���� �7ak�!x��E�wB\Ȅ���$TB�-?�8c�z=����ZD���B���A�+
~�Ϋ���`���
)�3'p�:�k����N��bݗ��u��}����KN:'Q� [��I��k۴�
�u������E|)Z��y+������"���W�q���6jl�7��=s�^H�ڠ#�r�T����B�{���:���H�z6tn���ED<dB�X����}ܹ���y���ku�bSP��.rE��_Z^5�G�x�̰��W	2����6i^!	�)[�(/�Ѹ���� t�t7�'�>��zIX��y5�[�uW��"��Wn��屁cw�C7�Q�7�%�~�������������� nA��g'�0�1�h�mS��3۷���.�A�N2l�՚�Fl��@f͎�W����8�u׺��q�f@��%�:���x\���d*}�o"�������SL���u��:9�­��:NL*C���ڮ;/������������[����B^����a�5�R	�.?���o|��^��b�$���h�m`a�*��H����PpX���ۦ�g���/�m���b<h(���B(�؆2x�輹^s<��u�'���ow)Tc2���;� ���I�y����K$��yEz��(�qY�5�11�oH�:�M��j�B��7�:�^��k+�g#ˇ)��,�b�Ȋ]��v�,~T�3��<��~��r�w���F\;��﫟�ܝ�1���!̫�S�J '���N��NO@��mZ�q��%r<�Oq(�&���fki<qdV�3�$C�V���5Ig���Y���Zu[�	ў���®rZ�wm���^�xe�����U�Ó�7��ԁn�)k�ѱ^؊y�vm�^1��)V\X��Es����)x�
RNcu7*��u����ő�'43I��b�ם2�}F��2W�y��@<�ic����>N��f�2Y]��Cz>B9��jP���bW�8��- H�D�
V��VS��G�[���~��s�/�����&�^��[�鈘���2��=�� Y_q��DY�Y���G6��Y���QM��9�(����'��9�xf/U� u�.�Rdk��m��k�R��,D&(���]�� H�[��s�
���O�__ �o����
�jxQ.��n�\��]z�s�@5�]t��ۉ����=�B�{���g5+:�<+�[�g�Z/���o�t�T��O�	S��Sǆ������j~K��G�W&[�.��q��#�^�ǩ|��OA�5�� �[G7�&�t�#�yW���Q"�/��{�0�龖���JS|d@F����4a%��|������zzA|q*D5wat{}~��?OωjA���-2h��6�� #�ɖ�׿��s�H��_�ϗ�g�B���/H�F�>'�I���$�i�@���7f�@��jED�~���"��1�qLX� ��R����~��<�7Wb�+� ٬u*��FLC)�?����r�� ���	E��x9��>�;f���a�\m?�$�a)����V�|�Ġ�C�/!��pC����X�B ��E�"��JQ>F��f3 ��cu�p%+~�2|p7`�J�ߜ��~a~�l��;�R�ul���6���	�{�D��[���|��-�Ue�rBAB�A����0خ�K1s��4$ ����@{�?= ��NŃ��~�'߃`���qa#X/tTJ��1aP*�JA�+b�m� B�	Tʪ��>O�[��_��S�<�b�Z������c�m��::���B�}`�ً�.1Pc�V��jd�b���$��|E� 1ټ]��J4ɺ�<4]�ܺ�	@
���@d�7�t�v�����^?O��tR�����ܔ��t����� 9Sxk*[h�����@6�ȣ%k�F���t���O����f�C#H��kSx6�����ܦ\�D�O�Ɲ�a��[�K^�D ��1$8��N��9�GZ�O��)��X�Y<b�V�ύz5�:�gb.j4�h�`�����`�d��"e�ɣX�7?�Y�D$A�CC�viN�2�n{B8�l����f��4���E*	h=���qQ�Z.�� �!'�w�/���F����~�Np���m�������"��w�_����╳*��*v�|=o_�=F#����0�a
8�4����i�K�é�1e^�4`�KxLj�so��K��J�ߖ��.���JǨ`�

��^fA�������7���-`�$� k�/�'�)�P� �bG��,��v-K��ϵ=ۄ(
o`�1q�GH�]����Gݔ�7�i˛\��
�
���GvE�s!jB����֤�v��ω�&�CL1�QH�F�_,d��e�΢�B���L�Kn�~ɐ��n�%��ZO	�9�)��]�S��r�J�n,E�J�@!�EI��	�h��K&�ԈY[^j7�ݛ��!��,s�4Qt3M�U*��:	�>dt��_��&����$-����셼2ߙK6i��6qk�h����\��_2n�Z3�<��+����'�Gh�����q���m�5)ȸv%y��$�Y�/-*�>��r;���N�K��zc�:�@Ǌg��&��ّ?ު�����7�f�*�fjܳ����y�璡�􏑙)!��h��l�AD2���k�w�&����1�/�P��aCd�� �@���<aG��	��?�9��B��>�ܢ�Ã[��a�9(�,���:P��9@��	��p�|�z͊76�҈$PD��>�B\�2:�w�ȵ��K���G�۞�!���_i5wRYԣ�m ŭ����o�B_l�5]�Ԑ� �&��m��3=�!VZ�cE�����ѓ�b�B�Y���${]#�w���"�e����F
K���JVPƺݴ2�an�J���1|ac
��0Y�H�H�����d�qx[%T5G�� sX[��[�*�(�hi��k[�;D�as��m�
M�j����?'��a"(�@�mTҘQ<�.��<;f4�g'?B������	'X	��!��Q� �4&�)(�O����٘c���!��*eJ�%��dkt#Y4}6�H+-qҺ��f��Ǟ~K4Uq0:���=�GrZ&C\Ȯ���K����u8	Zˮ���m�I�IU0$�N�^>\��aYrd��"6F���[�����9����ԛD{˟н�KcX���~�D��78{;�3�Q�&3_��0�w��cS�Q�Ĩ$^H�!�s0��%<�K����
�j.5���c�'����+��~����g�W*��o��,Eyq�@B����/�_I�Ӫ�i�g��c�����?l#ϐ&͈��뜕5fN���M�\�t;��z�E�ZrQ$�� *�؁�e��(�#�l�,Y��z��=^��4y�����3д�%�ޏE���8�"�I%6��}VQ�9�'_xh�� yD�Լ��O������d%<�:��Ơ�~��ď""u��X���*������>�DYW�GN�$
f����	�ec���;.v'��㺽����D��Р�A/t�W��&�M�#@�"R4FN����2�0�ra�p�j���Ѳ�I��0ʺ> k�;[ք��+0r�FT%(�v�-���;�q�AQ�� �!+�8*�"�6yj��:1&�K�,Bpq���J�FBM�o���δo���@p�1��i���<���DSB|L��8LR"�ABw��~]�J�vh��r�,�խ'���G�QQ��Y�%P�
����k��1��Z��"Q	�Nz>�.q���3FJ
ja2���B�(ѣ�=�$��s�0`di��pm���2��+����Y����2s�J˓vmH����U�aRR0L�Ӑ�Z;<}*�����^�ƍ�1�Uо��J�c�2H����F�Qc�|��} *~�P	%��Kt"5�+��I?�(�SP�0|�]q�>2j���&�|�!.w�� T
��B׷ �Ȅ	�S����"1�9����,3��{��>��	� �S��Mi�1�� L���7��5)P[M���9Gy�a{�B��¬Jh��Sy~�8+�͉-����>�@�!a�7#��[�0w�(��O%+�h<�)ƹ��ɠ2�mO�����v�(#��ݘ�?0m�+��|2c�dpt�y)�&�!H,�s �7@�hbz�¤��t�BF/Ch��F��po�����K�.o͎��I�_��p�BE4Nq���q������A9m?���H3����l��?%r��o�*J+N�*J�{�O�8��R�Z6�"	��͢�$G����d���+�kg�
\�
L�n���Fx`xt��+��ݯ�~��u�N>�.3hm�)�CY�M>O�]^�> ��r�)@�;,͗X�2ǡ*�Ƴ˸����rf
�&襳ן�����%+�˞�:k� �4�y����Z;�b�Ve�����sT���Ul��D�<E֑��M��1�_[[{\.��Y�'v�$
a,h�5#��5!�{q�dn�{c:�]V���i�|3�(AE�R9X6��ƀ��"Θ��6 -W�D�����%Խ�ݭ
�W��ȡD�"���KA����[�K����U#�/Ն��+��^��re���#d���ö�m��2����4�_6��_���
��Yp�{���	<��������Q�p3��������qF���9� ��k�:���y%�J��#`�:( l�'p��R��P���<��^�M��UK-t8d��C�����_DO�6�5-2!k�����p��0)5R�y�M|�hCu/Z��R��0*Gv���H�ly	C�3z�b��A	o�<�a� G�:�u�b��]��P`^��񋅚��%5G�9��?,� ��tD���mb|QvN�&J�p���:�5��I]Y:`�8�;�O��w_.�p/o�h;�:x�*s�U�^G�l�p���I<dd�?+���Z�x�mG}���;\۹����v�X>�׾/�k����@0��6F�m��g�/��u�mϼ����Ȳٲd�{�R��;�Y�@�M�$[�~� )
�<:,�d�d�<����^̀T�$�"��{�,D�,<�ijv���(cRm��3Ε5�H�fƔ�L��O8'����Z���S��rc�E�ͷ]��H5ܴj����F�mMހ+�Q���23�5�������'ohʆ�RP�6(�E	gB��B���M�s 4qH�T�`�D0`L�>	�
��IG B~���Qc�!@�v7 �
����!vb���_X��:M��w�����Z�4c��/QM�Wj =��ư�jA9U_f�@9Cy���I+���P`����|hc>(I$��Yoo�΀�l�x���I4� �싸a'~ȝ��'C$)<�Vѓ��%3W)^�i��b:�O��_i6���)���}p�Ņ|R���
oX��-���ޚgH��� ��pE�J��D�Y�@p�ƕ)�Q�XENl�h����rH�`k�5bR��9-E� Ր C2�8������/X�C��]L�
�PqF餝���k9ׁ{{��>Xα?{�׼��N��$>��� �Uz�+㯞b��Z���#+��]c�ˆ[�2��y��?;]����=4��ǯ���lIcS���?u�y���{��)x��S9F��ո�	���,9�^���`M�
 4_G�DLݴb�Ǌ�>�B�ۄ-GfyۇZQX�!J�B�Br��~�$�TF'�e��<\�p�T�7�<��%�y����0��J�tz�$��
�+?S/*x�f��ş�%�b�8CZz��;\:/7�Ql���]�X��l<��0��;q1��@X���f��Ƅy���X�f��1�'k���yXBm�6Qi+����#�Z�
���T������\Ï�~�8�*Ĉ�<���K�s���.̟vI��l���2=D���
Ka���V/�4�*/C�SgoT����7Q�C�]�;�ø��l�o�~*Xf�	�G�/���=�:��7��R�o��a�Q:��mc�x��f�'֪ż�����3H��Cu0��l�J��~9��A0�M���t�$z3�gG�P�(�� �ܻ�^��`:G���nژ7+k4���L��	�b{KT�j�F�� ,������ߥ	˫u%��Cy����:��Ǎ��'�c���c9eS.���	�?D����@�8X)(��R�,Ov��N���f�<0��
e�������F"�z{��Yp�>�F�H�������:b��5^�u�S����1.��!ڢ��G!a�9�B���N��A���j��&s��p�kM��X%x2K�ӯb*��W]P�c���d�� 3+��ε���u��8`��ວx[����b`�!DHQ�,=(����j+�6��������/o4���btF[�6�dm��
?9B >i#��;����|�psם�<~��Y�t��C�A�=B�o��/	j^�I��j�yN@�
zr�$U]���{�a���Rm���h�6���^�wϥ#�]�ؾ���@{=�=:$AA�q�'���(s��W�u�%8ǽD�1{��_�fl��9I��҈"�M�����jъ��6�p���{ n�[��h1"�z��$���67q�AU2\=m��(��,\q�����r�e���ܸ`]�-i+	�9u5$p�^'��9Ӣ�������ӡm��F�6t����v-���o�_�惇�����\�u@������m�D����W[�"�yد���{B��$�������mO%��l7�VW����BG"E�ΨCv{�h`Q���4_��wx����w����]�0�Ed�����M�oS[�%.j,�\.V=�8tz޷��k���*/����m3 8!��a` �xrN%n>�������R2�d"=�L}:ZGV� ��I�+����|�1S���O� �O��5N�|���r+tnFM�U}�:oPR�3Ћi���R���z!^������NWomh�����"D��(ԌKx����Gg�'đ����t�dH�F ��=�������״uk���J}��u6��Gb	ĕ�5���!�j�c���}��䶽[���fΞܭ��S���wG7O�(Θ�^4��m���	W	�ɭB��Cf�	�F���*j��";��ѻ
�������+y���sHF�kśH��xF(�Xh7b�^V?���-c��<Ʋ�9n�9��I��@���YO�1v/<��hQw����)��А�}���;|4>ɜA�������!'C-�9ݺh�7�O��j[�R�Mer�r{T���Φ@�M��Pi� A"'j��֝�f��F��k��I�;0HH-���%���O��*�04G����Ī:C���,E�34����y�.�0���ݦj�N����e8�3ނ��_i�UZ��V����7����A����2+p$)�H��v�S�����{�̸�[�U^w���^��yN�"e�m�áM�밦T�	� ������J��������pf�p|:�W9>�-�6��4n`�L �ޭ�$����'�1�L�)�8�un0Xނ�2Icⅱ���xLA���YA�zش���`�Ҹ-���߲���u�CV��SYcJ�����/h[�v|�n�4�1i2J��*��"/]�y�'<�qQb���ٵ�ZT�@M��G���&�}΍<7�sW���5M����']��{�>�U�E����n[�^j-��t��o�v�ww蔕X�\��_h�]�L�vⲾ�t�;�~,C|��b��=�qb��h̾�2&%�HD��9Lgc7A��Ch2�f�c?ݪ����dԸ�}�Fʄ��*A}��wIO�c��-Ěf�8�o�3I)��ʎ�(]��?o�5��+�~K[�Cx ���!n�h#^=Gu�����>s�n��I晃7`�!�]�$�{� Q��{���s�����t]=��A�P��?wZ�v:p��^نn,�����'���=����f��e��_/���#�F����^�C{!��6�6�۸%�^<n�l��aTv8��F!����}x�hva,��ЦZv�0�����ZK�*V���{&q��=k�b�?z<�����Yo��E�.��n�5��C �wwwwwwww��	�Npw�[~���{U�j�jwg����{�=�g��?�M��(0yK�1�Lv��*u��E6h��MuT�7�*Ȯ�|ȕ�Dl\�G���.w2���-S�q� ~Z����|Lgs��n�ŷ�:k/��G�{�6�	m݃�Kqs��K��I����$�O�l!�B#-��ă�j�y�bP_�a��.��K,��d/l�2��6�9�Qa�㉜��U���/h����l@�%�=*ZK��1W��V�ċ��2�����xE|5��<���)�-�\���=1��}���M�9���k�c���E)�7�V�U����N�9��Ӻ�_�l}H14�5�7�MU�=�8m� -�T�\�J�R�-tA�^�\-��%��..�/i$k�7[-��<�Q�
=�2G�8�����+�>�?�{|��(_l��xU�辆LR���W�����T���@�׏�X��0^��lg.x�����o[jp%uH��!��x$�S��1z�p>��ce�ٌ�k�`�B[r�8��Ka�6kFuD�����.��
e�*E˟TK�#l�D�[����R��Ƒr.� ��Qbv��*Q��P~@��>�d#��yj�~a!7���&�wܵ"�q�m�ڮ:Hg������N���m��'l��V���G#��%dR�呈�㠟�b8��`�̠�Z������Έ�9q�ݎeJX�Q�&�u����au�#t �>�P�ݫ�G�����ި�Hu�N��܄�]<�X�ӄ#�d�ڋ�����o�yL1�S�@Q`r=�3;,rH8!�� 8�,�ُ5�٬��}S���4�,u��^�]A%��<�x�캺N��x_���V����~S3�=X4�`�j{����'sm����m_1��H�UB��Բ]v)Q"��6���3rLr_��p[��p��������BK!�&�K�����wخ�Ko�ٜ���FW��(���"�b�s5�-֢�S��pc����r�r.���ɯzX�2���#��j��d���M#���"H�#��U�Fh�H�ZkJ�_��ߐ��c?�Q�;M��=�y����>"D>�y�� Q:J&�F�y`o uf�L������~>�~��Q 0����͎�_�+����bP�C6JI����T�q���n����u��q�m��j/�?��l5��	��H���a�z�)�q�Rf���iR/j1b�#��/�ׯ����C!��f}��4'��亵;���^d�/��%�X),8,����Z{f��IL���)�����Y���.r��[o�����>'1'&�0y�>���ꕍS<,���?�B�VyJXIe����U�`%69K���t���b�PluUsD�����	1!:���I��� ����_s�;m�3q���X��,"T_�.->`��^�v'���.��Vq������y@��y�0B�e%�A���X45&����iV~�g^R��WZ���t8),��$Ðӷ0ҽo~D�6"�����O�-q7LƓl�;��?f�c�ٝ�[]��[U%�W%y��U�� ��<{�V�ǣ�/J�!���.���|#����kp�rON�}��"3U�#�Ms���|�G�r%��\���	���Y����^P�G�%���y�|Ք/v_:��im���{�iV4].vZ˒_���yc�
�D�Zz3e�`�vY"�bʣ��9JB�E�<�H^�F��k����F��)�@E��]jf��(�+��58�'��'g�R��������Wヂ��?Fz.X-C���N�O�f�h�X��H��DS�y>��hbv?��8��2���g�i�o���)ے{�B5���ds�8 ���)�8b�\�U��|��a�J��7#\�I���C�1.@ߗi�M�뾬A�Y�׉�$�d˟�zܪ�Hߦ
EJ�rIa��J���b䎦�J��a �F��Z�ʪ�-�)d��5�(�W��JQ�P�͆���uC"���G!���{��E�f ��� v���X����і��8vU�m�u�Ʉ�󴡜�)���ΰ�Fm{BC��ܿ�e�?��%bSa���;��;r�ГqU8�� �2Վq$i%��qj0�<�@-5!��}��!�H��U,ۛ#�A�/ʛ�n1=.*����]��.�R�ٕ��H�v�@��b���#��� �����'v �%PCLk":O.�_�7!M�p
�(�h�s*��eH����p��Xi���D� �(�h��E������[R��=c���%�oPzb���b�9�K��L�d�-=�^����b��@E���T�ͨ������K������24�M��
-ǝ�,����o�B�.y�Kvv��8F!I���;�1���{��q�.�+��z��oBZg~���*\�ď��V�76�X3���#�צ�[���Y)+��"�Y�(̎����_�Q�u.��Q�b�:59�jM:f���#����0�����J_*
�xK� �$�`Ie�Qq����yV���f�"�#�0�b�#X���_���n���y�k�O��	�v]�V-��j�S�rf3`��R�ԚY �耱��BN\FR�D@ӎV��]V������ËVR�+�Wa#�Z�W�����v�
�g�3�Mi��%e�'� ��Pm��M���ۥ��������F�I_pI��~�evX�4x���I�ƾ��oK<�F8��Ҵ���������~�feb�
�0�s�I�Q"�}�x����e��T�'�wZ���~,����u��l}oh�>v��������2�bñ�G��{�acMu����ULw*z%l��bsd��� s4��7���ƥ�q�ُ�&�[{���^%-����������^��s�n/���.�$��b��%lG�?)sOh�*4�M|�N��#�KXJ\�8X�0��5��Ѕ=�{�]���"��nfJ4��� ��L�(��#D��9Hug���@(���jׯ녔�#q��v��HhM9n`i�����n����Oi�n�w��'ʛa�}3n��N" M(��3��6�L� =�P��9���n��n{�?�7�Ȓ�e�C���c���i���E:b���)�[�m[qVE�����cjd7�G4��?g�v����u��g�E�ƔV�A���>0���oT�=�_��|bc��@���&�ѹÍ)"N������7S�n:�;��M�ͯ�mndpWt�h���]f]�����
2�?W�^g��øT1V��τj��;��Hn
��Z�P�&��ݦ3�p�8��t2�5��M�haޅu�Rj��5Hy���.��^������h/��Q<�<��\�ԓ�D~�La�N�F�� �������vmK%����-mȞ�ŷ����8��^��GN�2ρO�2wV�O�4�qFH!]^�
@�83�@)�G8��8�K�9�̦��s�ӓc,�_h
Y&���P�=L���um�ZQ�lo79��|I�||!�QZ�T�9�,4�5јVl|��T�y&I=��|1k�%�ل0S�"c��~�+Ľ����|]@��+�N�ã�~�ӄh'����	{/�.���|tĎ<zJ��J�m^�R=���e�Q���z�fg�Bգ�:l���X@-��JP�t.�*>�8�����}��K�D�0�,m_��"����l ���9?|�'�9)�%.R?���˙�W0�P2 cb�%�dm0b��9�l���O��@�,L��%4Ɏ���J����\7�E�=(`v���lP��Wu�2�S�Y�Ğ�lֵ�8���:x�z������*��S<� ڱ��agb���Jv8��s��4��Q���6?"d].���F�����С�|�[�)��H ����r�����2D�>�FѰ���KU^��I��h_QRE�9oO��8:o�*l��ͭ�-.�w���9c@����RL,��.d��$h��J�X�na8�1�Z�9v0�^ى�?�T�;F[jc�l�i0q	��(4�3����ߣӸ}�J�y1>���W��.�����	�#^�����똉J5����&�4`���~�e<@[5PE:�	�^ǫ�~ŕ�c�?E���p'T����_Z�t�@��5(e�٬��JW�1pg���%�G�}h�-U�X���af��q�b���<�-���[�=$�
�,�����+��+�a��q��ޏ�g�;	�;&��d�_p�4tx���F���2ܘ]ʫL����}�wN�<Ԋ�]t6[y��Ȑ��9R>`�����7��H�d-����T6TǀҾ`�&�����|UKsy�7}�I�7����Y|5�{��9a�x�p���*ineu���׶1������#jT�������*~7~j���t>I���� Q��j���7��ō9J�u>"D
͇����0��� W����[*��߈B�+ ΢�hDx|��h�b/ڑH:�� �nCC( ]���8_A:sGH���q���X���l�Xo�����n�&�m��iL��ٺ1��'-"`.,�c!���D�w�����J�����D��ZE���(��N�*��Ǡ�,)GE��}��{/@�/x�\u��,-b�0�G��_�+�%��]�\7��a,<��e\�-�n����խ���o@�����J�滋H�"�	JD�M2��s��Jx��t�а�]�����$a����-֚R2ʲ��Ώm��i���-p�Y����O��24k���T)�5�U��L�^��-����E[/�W�&��T~�xI]�p7)Y�GBѲ(�o��)�I���^;U�[<��7���P�V?�Ŋ��%�i&�թ���Q��L[��d'���؜|�3�&�=�*�XMp�?;J�Mz�x�m�2��(cuz�جG#�@��f�R�\�%�қ+���-!��[��0�֎�y=y�j�=����>�;y|�v+���-v��{i9���j(�v9Trs�->v���V��q$�\���l�s1����IǇv��0s+�ϮW��S��R^�(Ix��L��m~㟹�%Ć�q�GH'�|0�6O�.��>�e%w
f2�*��K�X*��̮D,Q}��~V�5�����'��2TR���v!J��w�������7:�'=!e^�>^!}|�{�9W����JMa?nJS���P���1�l�s����wKo��UZG�G�=����\[l.-�7��M�q�e�xjj�o� �CiV҄<7�����ќ�K�,Z4K��K�ݶ���ވ�:Z�oNbS�^��#��-[q"�N<i�!b�UQ$���\c�۟�Cs�W!x(��G��U�)a2v��5�cԊ�c�6�I� O9�\�]�QEk��2'.�|��u��wP6a$ƅ8�EH�|^�f���_�g'���ie-��FTWĶ�_��Q��Ir;#�;1�~{A�6)H��%���/�bb9Iϙc�W��1_m*W0��a�&��t��S����Ҭ.C�6��)��oQ��+`�CDp�Np�c��̘�3�tI�gO\}�����q�{��l�]V����%sb��t04�X,
�&�,��ف�/&�i��e �f\�1"sЖ�Z��*l��-[��[�a���E���:�] gr'P��7":VD����?'��;c7<?�k��H�z����iP�J�(u+w.�5�w�6|���@��S_]���	�~�^�o���Ϛv#�kxk������%��A���ҳ�X�ɉ�kK�uGE0�U��~ǧIߚk�tU경����hh�l�a���B��sM�s�rp�e����� ����	D6�;|�yt�l�X��9�ǃ�dT��H1
Tk���F��m��	#{b�#�E9L�a���'����D�:��S,9קϱv�$K�|�V�q !�J�sN��S��%aD)!� B$-�|c�f�'��"x����d�y�\���#Y�����&{�*ӓi���wֆ��\��p	1,��Ѩ~��*n���ЛX�i��[��<ZD��g��iU�-��V�n�Z((Q�A�I�ۦ)i��Sk�N u�F�L�1���
��Tl��i{�|������Y!�;�7)��ӱҳ��4�S�(�+M�Nm-��*��_!�r�z�B�[y�C�2�\��{�#nM�qIv�1	��c����V��b�W�h�&�H-O⤯�3�N����d�PA����+��g���'</������B�P$-�̼�`�[B�0f~O�z�X��;=vKs���k��&�������A֕��*߻�;3�࿺?B�q:���i3��;)@�S�(��쀌�I%҉CE-W/U�����9L�=�'��pY-�����X�uQ$ѩU���E/�DQq�fW�M�m>b���)Jmgs?@��A-�o��
���l�j*�*]>�$eǂlu�ٵ��5�Z�e�n� �"����+{9F!��1g�{�F��
U��`��)�'��%M��#\�sk`�SĮ��}3���1{��&�^�`'y�J^MY��?
$G
�$�'�"b���ha��o�}=W���`�/޸�ӟ<Ae���me�����x$��h	h}m�\�z�;���u�nBCs��9�ޜ�6nU��)8U?�,f݋%���I����Q�8�y$�"i`�^ұ0��뚧^������Wpc�l��5#�&�6B���fղps���qpi�Y��pv���um	�MRF�*P��#�,!��L��GD �	�2�X��e��������o��"�_��J.��Ԓ�d9�I����B!4��qw;����o��ar��($�ĥ���LG��f��UJ�L��E���f�c��,���YrtZڮ_����F��^���B�)pw^�w��}G,:��PC�����m�P�rY�_:�%��*�Tz��e���R1
�R&�c&#�&
Pj7J|�=�,�ӛ����Xy��)3Hb�7d-߽JĹ:�ut��D���4��~��w3��[浻���3�$��bY�ܟ���H*�y���cdKS0~c��@v3��Z��d0p@`g�p�c�#qDSB;����Jk���K������ލĪIO��+�[��M�����E�=5]L�qO�f����v&���,��\&�����&^��"wk_�6/�����'��ݕWh����F�9ոq��qL�+���ܨy�ti���]�ᢐ�ow�2Q�}���t�襏�T�,��ދ"rz���g��{���B�΃�+C�5�,y���k0@0$.
��b�;�laS�M��//�|S]��&V���-�\	�
Ib��Q���"�wg|��x�z���H�w�Υ��;��KiN����������	��-���?���\,�č"j{sS-͝{���һc��q�� �)f��']��-g����(�O ��S/�f$»S,g	������FN���j���u���9W�7� �=hHͤǯ���m�� p�}���`B��W�'����b�t�_>�_�D!�Q����4��νkzI-�L��#�Z~�;)���q�
=��P���%N~R�3J�MU��٦��`q����j�<`
�M&�ȃD���Sk����"q���f���i��tv���s�(0ahG�,����1/�[�����:R�"�-�ʢזk/M�k�߸�ܭ�G�M���+O�3���$�zЕ�{a0�+9E�ύ%B>�~���..�B�%`/:A���M��+O��[5~�[�3��_�����BvOe��e��K"�"m��D⿳甏����5j��g�yƆbu{�����Z�X�=�X$}\�.�SQ-�����/7E���豨5�Y�%g`<�~�y��y��_"�k�P�<�@�p{<�'�m��(�����T��m؈!*6��1�s��U�Gߑ�{�������W�	�qDTf�,�eu�@�f�������R\�{<l�1�<�W}FN@N���D;x��b
���vޘ@#�֞G�s��p%��B�׏�uW7��B�����*�ƭ��KC�zeGТ�Ұ���۩�\�A�E&�)_2C0dKj�3��<��*Mʛ�2ul����gJ&��b���o��֩��:�.x��!rq��:?�+��ä��\̔��ܯvɒN]��Lǝ����9Y  Z1Ls*2�m�)�J�{7�|����~����f#��A}�������nh葅*:<�Q<�g����3��j�v�0�ߞ���_-o������t1��P5fW�Q#08�y�ں�����'�����b%|�dz���-]���A��ҳSgɪ���x��G����]�=��>#�n������z�Y�$�$f2jYؼdTk�j�Ȩۺ�>��H��Y�z}�'cv��S���Cbr�0c]��zb�c�S{}�Jq��R���8s~'�rg���z�_B�_&eϚ(�&����k�Z(�'�L���e�yND��r#sf"!���.9´�#������N�l�W��0�>j*Z̙��l���|$c��.��<	#�K�t�%�]�w�W��d6\���E�!h��cQ���+TǱ��J��)g*�AO#߫)@�F����#j��Dv��8�1�#�������
���������q ���C���{� �Ĝ���mT��N)�bN� � u��T$h�TA��!�O0�>;
m�l=�+9o��i	$ĺ���L�9X��]C���!#��U�Ow`���_��u�1I<B�G'h����j��ȇ����������;�y�/�c��M4����D���Wr-g���TOT��x�Wqɑ��	{O(A��a3�\�to���F�l�d�)`�/���9$�1Sy � mؾ4iYzѼ� 2�N-U ��v
�� ���O���w�G��O:,\��z�|���������=�U��W�K�?^�N�9��&���
̹��D%�.ѐ����-���r/��8��0R�e�����3�t=}98)�PY]tb�1��K�U���&�-F��:YAyg&���'�?_Y�[�C2-;:$K�J)~`�SN��8n���Mi	���%	cA�����
�y���?W�B�e>Uf�t�({�����d_�\ŬI+#+1;��fD6��Y�Vj#��Y�L,Cf��/YCoȃ��P�5�AJď���<a�X�����Ȭ���SN�L��z�1r��&�p�3d.dm�;�e�_z)���?���<�S�嗕�b�/^��A�geM�R$D����1�Ox�!��3�#pKv����aT&;��U�c)޿��8/�����%%�h��|�j�i"��@#����槟�ŭ�
	ꏜ�^{BHaRԸ��r�ɼ�{qq��hF��/r>��~���.��G��f�G���L�LYk1�qY��g�J�LS��u��P�!pL��_{�Ĺ�P�ٵx����nL�n#�z?��q�[/�Z���*�����"�c�����e�]�{�2�ȂPəE0����,5/ϲa��җڌ8U�L��6��W�2eM����pG�3#�5�|X��+���"O#DôZ��5��pk�(�0�e�����0��M&(j�J��䪟�k?�����dْ�ēz����~QT�͇�������P�]R)�;�P.�nν�ϻ.��Τ�{���0v���B����¦�m�a;#��T��=���͗�&+���ݷ���w�8Ʋ�<<מ��41+��+{)��z*~��ASJ2䍄KV���JJ��&m*�9�ЂT
8  U��ͩAEh|�e�Pj>����OW��9�T�}@�\��9,�t40ș�}g~�p�K��*hV�)�$)���>>��DC���E�@�x�gE��1�X��s���i�E��ؔ�6˻�Iv�l&��r�����& ���筇j�k5�Ъ':����-��o�P�g�����c���e:/;Cr<�#'����w�=��H��0�L�hJ�~ ~���Qo�)�Ջ؁����?oMtDx�1���g..�;G�z1�R*>x;�u}�>����歐"ah��[��x%@a����|�������(Ll ���/���1izI�!�4�:(���v0�h�����ï;wU��{�6|���{�Qq׫X�q��Z�m3M��1k������P[p>�����V'hP��(p5��Q���,�� %��+����&eg^��������L�Gw���X\
��)�q��r�O�$Vo�������'�4�7˂e_�ּ�_��2k��-�1"D\�)���
��X���aq+m�(��u+]���G1�*g[�k5W��^�������;X�ͭ\	I�@"d#Z��4��K3��
��Q���U./��Iw�e|z�eSl;\������x�:K���J~Td��>���r�uPuh��ד�_1�#�ƨ����kbJ���p���" ��t�PW���u*�&�I��4���E~z?'Kǉ+_>�߭x�P)R$b<� I�
Il�´]�������p�:�[���������PM9*a;����z�PRD��>�਀����=���p\��v���N^
LxLx,5�����G ?=?1��$SK� �ګ]��*F�l����ϊ����ˡ���]���������~9o!X���Je���-��M40ޑ��D~  �VLPL؊���WH��i�F��hX�O�=�K/ �A�%��Ȫz6^�R��q`0�bd��ۥ��x��b� ��Q���<�ta�N�qX���H<�E�-�t��L������F�J�}�<�0���%�v�8��v<ѩ�"��eZ���@C.O�������`6d�[�� ( .�����F��%��'ؒ����Y��cs�m#EH�/�^G��kik���ʡV�1HmZ2����k�����^9��x1�"�˺�~���V�Um��ڢfG�
�A��(�D�__B]�U��u� X/��������nb̌��H�T�P4�+Ѽɔ
�e����fz�-C�K��WSx�qh�儚��m��0�\#c�&:cZav���ƑL�eX��R�_8�Zk(�(�MŪ��6�#�q-��~�����	��Z���c�MA�y�E3����E�V,[��(s_Sf�ik�2�>��SA����cg���E���ݍIU4������e���\� ��_�Ѡ3��������%S��T<�(A��e�����rG����J����i��[f�v�0:�D�kE2���m�F�B�m�K� K����B�x��x��@�7�g���ŀh �2��πx�`9b�	3$3#!A�xi���Q�f�'�@r%����u�#Z�cƔSH�n�"����#{��O��CVB)=`d��H�U
���d�����&i�����W��F�Hhp���)}�+���B����9J�������Y�>z$�;���IH�(��tc���^ϊ(��k�A�[5��:�b��)������ ��mPI�g!����i�	� Ɓﭡuud7X����Q�Q6l���� &P0D��k�1Q�1�ݠ��#U���/��	W�4�~���|����������#0��]I}���~22�8ZN2��2#q��|�P9	��=
�H/����C]s���O��WD�;��B��f#�ϻy�ʳ�r?\�ӻx�y���&���pX�#���ٮl/�cW�O�?xF�֎�֮l�+I�+ǁ5l�~C��|׆�zX�jF�CՅ���?r�?��$�%��[%�ȋ@�zbB^�L�����(�$��͛ޢݪw�@�:߅��Txa�p�����p�a�XwJ�R�':��!����Sb����P�|h/n�?)�5Cd�,��Mb�ߠ}fŊ,�W���H�|+�0�^�:�;G������Waq�~�_��/4)��E���Ç�Aq��5+Uho33��$lt����S��|qFJ������9����[O�g
T}��8h��Q9�P�/Q!�Z�י,ĥ�߆��A���q��9��cbs��#U�h"���D�5�����季47i�Pf��ry�L��-���y��u�gcN ��R-��<2�����-+�K.
�������m�p48(��bwkw��/E
�b�+�p�tL����,uP�@�G}�LfE�"(ѽ��9dm�7;�s=�bD?�nD��f���6�L~j��n���{�׫᧸�.�uю�`�xΨ���`oE[$�����v�ؓ���r��^�ʙ����<ݩ�1X�ʐۇ�ё1��a��M�r�)��=�7���eOj�_�n�[qVcR���k�"�'RS͆^t�q���6������F5��Ϯ���z�X���f��l���e�f�:�>|<�?��{�|��k
 ]#�a9��F����GBKb+��h��L9��x��K�Cػ�������2�<8Ć��y��u�^�~�7���5q�@w�G�d����;o���oy�K.��1�}X��QTh��Jܲ���j�H�M���7���-$|��\>O]��(���ܽ�7�2;����y�<>(m�w��l�� &��X��V�$�"i�c��	��K�Pt8��5��5���"!s���Aqpb`�}r��;@���Y@����T�P��ϡ�j`[C�_R~�4aG܃���n$�/��������/U����W�߆=%�-�B>O]�����<ޠ0�[�.X$z�`���>�XXx�Do���0����sx��T����zO��f!�/�VoC�QZ'>��5�;��p�����٠3*L���Y�Oɛ�/h=�(b�GHl"0�,x�,�	$o7�AHm��,kM9Tcc'6*�V��Q����LM��u�X���t�p1��x��s���"�Q�k#��� tRI��.5=��D���"*�G���n�ϣ�DC2���WR�k%R9A"��w��

&TM�0���kZ�g�#Cm0<ZJ9�䢳�j� �:1����;���n��GJ톌�hS�	A��/�(i!Ԭj
Ʒ�XQ�n��y������\	�"rҐ�����U�l�@@�耔?�U���$�����?뚌K��,��7��#�<Ba�M���c�������	v�j��Bl�����������v%5<b=r�j����ك��3�Ա@�b������inQ"a#נ�a�$��.\_8b�n0��ē��+� ����"�Y&�
V
�n�x�]`��?-�@-b০ޭ௠�h��s�&Ip�?MP�YU��_�U�>�D�W�'�^[͸��J�7�� �\B�!�����48�9��̥�F�:f	t��vZ�]�o��q�a
������՚ax2����԰n}X���Y��^�A���&5�M�
�X�O=^5��ضN���*W� e�����4u��Ll����F����n�i���h������0[H�]	?G����@.j�Ttàı�+d��rO��� �c�-��OF�+�T��ϣ�9X�
3��Թ6J�軱�i&C�G�Eώݘ��g��I��\J+(�z5l�s¹3q���2S�b����ҹ;\���F5�:oF���&��0��!rWf��5��Ħ+J3� "�{��P���r�|�Ⱥ��B���yz��%���LF���o�`��M�T͢DE�zp%�
x��[~����$��i\f��1�ǖ!B+!|��_�(-��.a�O�~҂I'��Q+gWF[�ȉ8h���~��{��;-���9=ul���W��N�v+�>�z���*�R9AZ�=��x�'����*{�[��k�䷴�� �bu!sZUC-�a��g:p�:�+T������=�Q�v�B��@�S�t��R�ڄF��^橜�e(��݂)��1�����t׮qiΟUmڷX���=�Nz�$H�9t���1X�B�X>�P}�?��d\��	ʎy��xZA���1M�%��U)�ک�[�U섎�@gB�Y(d�7}�����[Hn��lPQ��2vvĘx��&�i��{+�X�"�'�����=2
�i�`�U,b�gf����G�l��"�#����xI�;��鈸��A�,5;@F����*�P�m��&���������V�k~��K�- ��p���x�n:�>t)� x��M3�)�M�l8�-����KG����8�`UI?���`s�F�p�2�}Z�����O�Kc�f�
�!pӪD%���׷�H�
�8}�Q/�`��>z;C���49fjEPo���X�Dr��;�5���^�[� A67�>X�R�ny�7i<��PI˞S��xMx��n�X�_��O4�d׽�0[Pr�eT��⽬�k3<nvGV�P�^.�/{5^�r[f̉�6�y��y��E�YE�G���*���Ur��%���`��Y
�Ʃ�@�����F1n5�}�z]��<.�W��D,J�d銛a݇�Toud���:D��Y�$��6�+i*$�C��`�S�ws�c'�]!L����qZ0<��Ȃ�u�Nw<�����D��Uo9�i��ş"R�!��,;�6�\(Ճ>�X�>�"\祫=�Ǿ2���`����_i��S̹�1� :#��j\�����[�'��f���ن�V㴴"veў135=���	����ɧ��� M��`���c�5|J��i���'E�)27�J�㯐$b�)��B&)U!���f��A�m�4�!b͆�qi��}�����J��9O���n�8��
�tF^PG���x�\�x�[c�v�RP"?SJы"��q�r����$��Y�l�(�-�P�J1��^	CM}h�T0��	�P�Cj]�P���C}a&��l���Rگh�����@H�.ޮ<ֹuSC�˻Y��h�Ш��R���.���=�C�X�;�J%V�ik�W���z�m�z1$ވФF^�7^�'ۂ�1����j�B�tJ`q~g!t )c!�B��|�-�k!�Q��O\�'��72L+�|��[9�VX�7ڤ]<e?K/��@/W�Z ���d_-Du?Z�s�S2�&:�#�$������tJCe��U��M��;��F��x�jdwv��ѐ�8��7�
�����1��9�-����"ɅR���48k�nն-��\d�p�=��zd)�hk����ۧ��+ �mT�v>�w�t��7=z�ʁ� H3���F�K�#L����@l�[Q�����6�2d<���'D�T�F���-mV+�#�&��0K�R���k	׬��P[f�_AnWL�ˑ�U*�u����$�zfz��F�Ah���B�Ǌ7x����ݰ"�ne��u5�B<7�++�����20ŎW�6�<����ܑuk�����\�@�B�)+���k���M���J�\KFg�"T�"�E� h%�#�T�  ����x�B�,\�b(g;���}]�@~ݍa��V���$��]�+9��FM.I���7��3Lp�e��sfn϶���bs�+������X�4�y��� ������8�����"�$�	f��ri�3������MǗ�W*����P��'R�t"V>�!H��.�҃e��8���ܳs1�� �뚋��k�6'}b̧���3�!.ko/DK�[Q#g7��e�
�E	�zzh~�p��7LP���-fv4��?�L������5��zw������Lӂv�~�F�:xe�~��;R�r��|<7Dת.c�~(r�h�r.� 1O�$� 3u�fj����(3m����N�>�l�|o�)]!�K�r��?�F�ڋM�~��u�������K�$��8A���F�ۂB����E����z���%:|���Tcnt�Ve��=�)[�p(���O>2�W���u�m��Nt�>>H����_C
�k�S������I�/��l�4B(������Q�lcNx���#S6A�s�d�m��6j�-�-,�C�7�Mr�x�61/x ��QPR�L�㱥��;�m��(=���
�#���ǥ%Q>���/|��O�,����F����\T��L���k~j���@�����u�.�"	������G���Qͭ��a��:��e���>�6���m�NU�1���a/�����d�-�p�ȟ�t$*x�hgl���{X��[7#�3K�*�~��Y��RN�7*+�	���J����L�������Ȏ�rO>x"�.[M_�	_���/��SD3���/�K�+Q)�РK]���ճʈ� S�K�gf�܀+�D�k�y8x���o@ݬ�	(����|�#� w�8
l>��������3
���f&����Z)�ϲ�"a��V�����' �=��e c�8����]������0�O�h��y�"�������W3M�A��\0)k�ET3�q�0���>ҳ�=FY~>�����:9�_t] �;�ne��O��/�X��R: ����uЛ�Б��ۨ
��na��y�&�{�RO�]��p�>��[
�R>�����I�d:�H�N�1�ż��՚ghM��h��_""���<��lHaoh�/RW�;%��Q���g�J�r�
�F6�1�9x�m�����+���0ww	��������5��;!�����n�/�n�{ﮮj�v�gG���z��y�?(訩P]�Se�[�P�x����8�>��R
e��c^MI��T���7�#�ʌt4���h�#U��NKv%�9L�U�.��9�U����6��V�B\�ِ��H��b��}����"y)��tϢ����m�[��^L~ng�p���;D��|�fYg�՚�Z; -<O2.���{�;�� >���Sr�$f�X�db�ߧ��sP4�AF(8EH�v�ӧ�%��&T*T�u㋐R�tI�=�����U�|L�f��]xL�.mL){Bh���$�-)�{���ǩ�M�++�M��d��G��ik����@%߬5B���Tk��#l��$
y��f� �����*~�~	�h�*=Y��fܢٴg���ǐy�Cذ�	gT�F������~*gC 54�C�/��$6���y3�^yG���>L��C_���W#2�#���8"�V����z��hm&7��sD����T� �e��Js�@��OC�ov�$t�)� ��*�@�Xտ�$�����%�Ù	`<g,Ql,�����S�2h�U�|���e��Z2]C;���s��N�7ҕc�~�Q:B�$C[���F�dn@L����X��/��;i����%��~l�*���L�G����k�
ޕ�F'�)�1cD�9'Ș���f$���F��ؤ�W�_�c�>oz�$񾅴�E��0�����*�7Su���G�]��3(�U
��'�@x�*-�^чY�ʎg�!�Rѹ|gCĞ8�̈ޣA�
����o�J�%�)~�R�x�%I/��̷�I1C<��20�kg��Ӵ�l��i�d��CM�3�_�D�<�|e��O�kII�_%�j�^7���L��ߐ7�T����B�є�D�C�|�`(����e�B��8�-���F�G>��2�E�	���K���C
�t���$C��;�5�uQ�!.rX�W}�҃�YU��8ԳZ�&�{��ږ��x�v�Nɬ�;S@�G�P���%���d���x�|g�}�t�a�OWC!�R���~V+�P����o�HkbX-\5��՘�H4�%e񵓥����~�����/nO�[f9�n���	�,	�x��r��Qgְ	�(�pH��$�5n�>(�}��'7Ϭ�{q~�솳Xı���!�\�����.$h>� X��S;ђ�o�~����a:��c��pzT��榳����\|U0L;���L�pK��%���s��.���v:k6�ٱ�R���T���3���Lsь���K�o�9�����s7�\~�C�f�*�h"m�QQFK1����V�u�0�,�#��Nvc}���xC�9P��C�_8����^�&<`L��E5�ٽ}�޾%�_zJ��dP�7��C�U{s�SP� -�e�l�hG��p�T-�Q��:��tw��d�f��j�\�"L�����'�е�d�з���J�P�B-�Y�Uh~-�� ?nrN\���8�u3�7�z�^jԷ?�_i�uJ�~ū�)�����nL�]����`�:`��|�թ��+�l����+��k��'�R�h.��;���**#�0��,�D���78�)��%F���EV�*����C5@����P]s���	I��Q���o�i!=�A3p�h��I���
e�߰R�y�oR���KF�^R���1�����y���� ۛ�I�(Π�W���8�#m)K����ۃ���x���=-������nS�8��ܟZ�&�D��4{d����;:?d�T��z�����k��I��Z�����an:��ԌP�����7�g�c�fE�5�[���M#G��D�<U�����S��0D��ԁw��+TDi���)6;CF��5y&Fzc	2�sr1R�p&�����鮆R60��T��s��\����|�~��������U��cs�ϝ�>]��ރ=.�i�g	���n�x_���BI�L���IoƔ�C�^������RVDY���ܞ�����5�^�
ˏT�|��5��T
�Ԃ���TTV��t�G�)���6>e�|g���	I8�Fm���S���^[�n2@��ݎ���R/O�+$��nn�-�@,	�����}���`n���4F߅Rw�� |�� ���X%�R~�T%nLO6	��4�df�w��[��,!�[Du��UŬn��!-�����u�N��ςz�m��\9����wh�`i���,�Ҁ[jz�3h�rLJ�0vۄ����[h�+��FE��}A{Rp;����~f<t��	��Qmk�Ty��	����ַ=��AcB�%�#�c�8
��?�m�v�	�N�VT�3��C��}��Yẜ} 
��(J 0�C$�V��+	\�w�%�'T����l<��m��G�#�Y�.#>a�X5��q$��E�����D���`�{+�#,��:yi�8�=)��嬿V޺~��m�������:b�E�$�*�Hۆw�Z)�n��t��� �p�!��q�B�"��椴�X�Bx/Sx#��4x���4������*�ɟ�`@;�$� �zU��M�(rtd
��u}��d��/�J�3Oy��T��s����l>|p*䣆j2E����"p�N$��H\h��F��?֯,ܘ��P���+R��*w�P%��o�I�i,׎��a�ƫ�������$	�����.�RǦ���>���,�D҄&���G��k���w #�
á|�6�µ� |R�._@ _�FV�>>W#/������_B>n�S���J*fk$p���|�K�j(��8�Xǖa�x��q��eG1}�3
�//I�:;��	\����8Zr�����rE/�t!@fu �^������?-�q�I�F��s
[~�����CS,&�����&�0fp���ٯz��H������=o�;��vgUř�WĂh�@�5q޻�0j�d`�O���ձu1����e�y��!��dZ��`~Ÿ����C'�MR�t`��#h�#.G����v����*?/�����^�
�N�^8��O�2������&��6d ��w�m�LK�c����pS��Z�ڨՌ+KP�`p���=�ТY ���1W��9V��?\�����\�R�\�V�s���-��av:}�*�����[�s9����EQ֏>�/�	?��f�̻[��	�!%MW��xm�d"�Q�SJ��� i(�A��~�Oo���#s�&A���|�ЁDϥs0>}��r!�*��D4˗5(W��|��W>�G�ợ4��f4/��e�s��l�I��H���]�t,ymo�~Տ�Nr��t�=�Z`n8�4���k�L��Y����������{vN8?�0�z"�G�W���`<����5���>�,.��(d[3B�:K �;E���`C��hO��,�$�J��"%���X��q��"�.v1���iP���Oc|�C���.�+�m�c��|ٰ`k��ƈ�k$�� tC�e6|nի��4L�'>�t�e�-�$z~���;���+�ֽ��Rm���ZZ�w ���JM`��&�Q��h@�U)%���yj��0�G��n��eo�~��m qE;C�;# ���/���B=�,"�
'@�%��G@{���:�J�:7��E��=���Ly��s�ߏ��\!�~sv����F@"թ���5���"�I�|����n)�&�ϡ���s��9Tb��OPվ�s��"s^�5�%�A����D��p�FY��O���Ѱ2�rI���h>������s���]o�TR�߽�u��z��������t���"��ڱ����?�p�a�fT���=�r�&Y�ݑ!����S�G���bw���k���(o��x
�d<�+&m�D�"�ȰPK�{��p��ѡ��M��S@�q}�=h�ׄ�y>L�����깴u����A*W����0K�M?�/ j��m��{T���>xVf}m���rh���\��\�U��pl�XE.�l�H6�Js_����>������8���iX6 -z�˴��n����MH7b�����7[8��M���K"�`����d is0I�hQ-����,؋�Z�:c�ݛbqk� ��{�|�����e�������M.s�����	��3�ϥ�� 	hW��9с ��k�=�|8����ȡ�X���Ĉ�s��wmQ�&R���[�^t��7��m�%�u>-iӌ��V?�`�����c���ܴ��x���OtZ�@n6ȁ��o���ra$����\|���)���s@����)����/�$�3�*	��f�9��uz��
����n(WG
0Fj}��[@<&���q��lq�L��[{I	�ޝ+���w<�����KK�Ʌʱ�ރ����E�7�ű�&	���%��-lHZ<����t������PX�mݤ�����d$D}K��5�%�+�L����Wk��mG� ���]�)��G������m��n6�L�f��[IX�}T	�]Hl��(S�����:=gư��I��۸�N�'��]�!e�pG=��Iq]����C��bܓ��U�����2����+m��{�`jq�h�FYv��Ajn.|��B�"0^�.�!;�<)��\3ˀ���.Kjr"�gCu�md;]i4m�?!/�ܾ�$��N7�X��1���CDOBM�8k�A�e2-6k��&�{˓��Om��My�ywvv�����H�|�)��TgF%�'��=k��=��ïA�`�KQ�ZT7q\2vk��U[�!��7O?��]"��a�n-��:�#R��������)�x0�3_f��
�D
��a��NoM����wx^���S1� �߲�.9��_��MK�v�aJ�x��d�
�,Y�X�ȫ��N�=�]�7E�3�E�l}J\MCV�#�b�>��=�CM7���c���t��A#/3W
����M0�[VP.�{����9�� ���Ck�O���h������OvEߘ�̷��&�I����E4WcY+���s��.7]>t<N@ J���g�z���Fce���)||�.��Q�5�,��*��$�C�v�Z 範g��d�ໂ�z�-Ԯ�#�a�T,�h�[�*K�P=��C<o����u��B,��	�N�����k��6�z8z�y�L�ʏ��ټ��S��('u������hؓJ�oع�ȅ!ӑ$�O��JM��P��!�Y3��Ƚ�3����ɟ{�,9�{��Z�����������d���:�Rˠ��%�e�bg��uD\𖾇��gf��8���
�[qI��d؜�P�.����4'H��P.�Q%|t?��"�w;��Ҽ5�D�l�&�Sh�J��Q��F��~L?�ȉm�s!�A��Z)�޹E��{ۇ�G���8������{���J�� ���E�#�������Rb+�4`L6�G�|��F�K?��r�g��IWйH^�q-Mn�s=u�۔�d���3�&P)�t����O������x����I�g%~6���Y=������5�9z1>b��O�G�w?Q�|�LP��l��U֢|��#Tc#N:#C�|�v�\>>�Dk�W_7�&P�+����^�>y�ݳ���W'�Dfh@5�³mнVe����[K��B�6���]���u�JJ�B�:9e�q7����/��3*�r���8��B�GjwP�G�U�)��ſ,��:W�;��qaݩ8`�������%WQp�])���Hʼ���G:� ���ViN��S�D+��b�6�?�a���3?]*�r>h��<��������݁nX��"r�*���Ɩ��˕|� Z�A o:�?�x����>2�~���l�#ξ3y(��3�V��� �Ԣ�
���7�Ᏹ̙8��L����徾��q�U�s>�p-�٥{,�˔x��g�Z���]բ���/���,���՝���qsu��`BHþ����5�[�ԅ�������|�A$�a6�$fB���Q���5�x;�F��G���c�B�
��6";ĺ���
��oW/h�3�x�K`����\c�Bם�ul�s�)﫠et���[�U䌄������&�܌n̯g���(`�E��rqqI%ѵ�n��G��$p������Ͷԩ�\ �e���R74990�؂;�+ֺ�����W�3h��էBO;/Jb��<��������[�j���刍3�cM���B���⺫�Z�|�s�7��}�[���Sjf!���sy��`\X�ɾ�~^�k�VeI;5�=R%���V �g�#Tk���C/��i��!KL6����ˤ�h-�)cv�5�g�QB9uz�>�0D4к������U����u�aA�ns�KE���Y-���:P�I];�����@���/t�=.�r�6�ʧlj/}�'_1�
���P��7� ���S�l�����r���$!d��tpXr"�Z]�]��^N�(@���9��t[�Qvz@��fD|���$����Q��{`Ne��k^l���`YJ�=s�%oqg����������៾��;��^s��ȥϴL;�e1L��(�1|��{���w9!n'h��'�]3h�]���
�
:NЋ������|�A��wd�(��T9�c�s��*�M�sd�����7�To�a�.Au���H�gZ <]��ĭqǍ���C+����廁ҷ?�ڪ���&�bp�)~��2�/ʸ��45�e�Ҩe�h����3߹�<O�`�F��ߑU��0Կ�z�q�I�ND��w�xq����PP4�d�n�]�<,���xI�:)I�ވt�|�o�7P��?H���cסMA�t%C*U&�m�����J�i�ONI���9�%�S�����y�H�֮v�IU����bEq'��<�"CKh�,��IM�<��NȆ�h1@p�8�D��t& tlg=<�X��ИKԡC��;���{p��!����Gڎ�������o������3��j+B�����۰�f3snbxU�|����3p���}�
ɓ%�I��n�N������M�&�8�ZP��eԸeذylKM��.B�"@���*'��M�
��=�CR��&�C��CY��5��M�n�
�.}� T�<!��s��(�G�f8�+���S�'e~���$�-j�yk4}s(�
��F�:���{�!ʫ+�D*6g����PTs1�5��l�uR�&O������d5�9�И�=rũɱg�)B���ir�{8#q�����3CX�{�f��M%�x`�'�BP� �K���lI�����9����_���9� SG�;���0O�<�z>�f� �]������D
�f+�����wEy�ǔ���-��'0��w���,�ʌ޿1�ډ�� ��d�	L��䧘],��|�'P����S)Q�;mTq�О�H��.�Y������Y�/�������� òu���j�b!P�4,�6c<ܩIs�6����x�ݹ1��ڎ��J�,� ��%���18t��E�&l�4<E����F�[�5^ٟmvf�2��˷p� � ���<��P靯���˸dG�>\w,�F������W�^E���Jx;��=���/&u�7u��r���A���|���ɼ�0��1���r4<�w����ƪ���YE����z��S}HYY �҈T��Z���/�:�E̰qI����:���h��;��OƗi��Y9t�w_ �|U����x�]�;�Q��<�?��<a�C�-����Ҟ���E�X�|Ę�{�rL����ƽ�����'��$v�I���l%!JU��G,F.�"�|P��i7<���G91�����-|Q��:�W����)`��2��ǔ������^�t�O+�X���xzY��1ҋ$�|ْ|�>3m��0����/��^��6	�(��V6A����z���������g�v0xY�X8
Z$X���t���Di�1�.�2�[ק�ݧlT��\���G;�s$ǋ�S	Q��2��H�	���Y΢e��}W=U�ߓĹ�	�oN4+��=Ĕ��}�Y��J�T궴%�3���x��t���]�27OQ�>�*�7�`0)ǽ���Jo:s���K��@��W�f�x��y�z90$�����ǿ�Ym�Z
e~�§�$�l$��\�
�lb�o-�l;w]>D�a&iMM��r�^�l^�	N���>.5�|H��o�.�� ѥ�}*����.������ɚ���-�o�]��&6�`�1��-��P]��k��.s�������P<�
���~��:O�6������.�<���?8�@W��@dg���n�F�{vl�b�d(�6l[�h}�8#�O@K��� e�'���$����-��M�(nv�b�"���R�[�~���gCSQ�Qsr��� QpL�S*H"�5�g�)����~����wlHO0�1�yZ��"F���@�'�o��9�]�o��Ij<�@?�Xyd�A�z�HF����C�����V�"�tч�ͬ���)s�n�g��6@9���}����1��	(�-] /�Nk
��߯n�?�!��8QL���\�dG��xx�z;��L{��aS$���|�2_֛޽��N_��/��5�o|=^7iz�8_1����f� w�#4��x39���z�)a�ڿ�$�t��wH��ƈ�7*�V�(�.Nn����Q���b[���ӿ�w"��.�vP�w���]���2� �v���\�V-*,e�=���]�s� ��8��;�#|�fߢ��t��;N[�C�ݐ�ܠ0?`�Ƌ0�wQ����"�M�<K~ޝ�}��"kn:�*-�'�����Z��5�����/���;�S��u�v\�my�!h���H�Ò?S��m��
1�����-%��v��>���0������q��֖0�Y�X.��f�{���N�%�@���"0n��_��$�V7�>��&����u3P�&�w9�I9�{�c\>�s��4O�·C��W��Fe�U!�V����Ȫ�av���GHN��T~�����g�����R��V��� ﯚN֝�v�7�</�=#�!$�[X���?�����ޘ�<`CJ��ú#�31Z�nD4�a���1�����*h�>^O��כ���K��^�V~�;�0�c 1`�w�Phi�%԰�V絹풦�����K��E�1�H�����W���nHJFUTk����0t}�Jn�EѸ�U��)�M4>�x@{` g4��%��xC����R��R��d!�t��c��d��["ᷱ�HK�޴ o�KM�uqK�� ������b��)�5��f{yK�b�K�g�j�����^��A�c��ȍ�C� H@���F���jѡ�VԀ��R���_����]�U�l��)��������dN�|���C�?�+G��9�W��61�jn�����V1�Z�G�ձ���hE	>C�ӫ�e2N���rw�o��s�RVQO���z�'w�]���Bk�{�?��=�Q=;����?��(Д7]n=H%�9ONϒ2��a�� �b� ��8Zi�p��^�v����#m�8�E.m)�Q�b2g��~S����>��evp�A_Z����r)Ó�?3z6�me���O��z��xn0|�*dE߇����0�r_��%�z<����#u!�~�;ۜ^�JF��X�"ҩ�v��ޣda��]��l����8t���F"�V�Zl�M;C&�9���{E���O��vjs����2L � ��7�v<��>��e��������9ݥ��+q&\�����V���7r�%�-�ѥ����ԉ��X�i���?Ü��.K�����J���ѯ\�Z4U���l�$P ֳ��O�O2�#�r9۬f�6��;>�xH=j�DR�)�h}MZ��C^�u�k�8��,l�����;Sߌ�����{�䟋EK�,�[	OSaGN_������TR�����S�@��6��Ow{��
��<�%c�<ޕ��|M;p#Ƥb���#�V� �,����+L�P嫯s��k��1a=,�JNcP>]��\'�.�A1J��u,���������/ˊ��q���o�.*/�co��[�Y�R��-�&�Vq�*h8�dcW����#Y��tX�ۂ�Jo�z��=�0�e
*&�S!�q�����$������k��4=|_��8T�c»����a䤒[W��Th=�}��;a�U$򡚘~N�HtRi�6m��ᬽ^c�z5g'?&f閑�OV���1�� 4mZ�+�2z%#B�BE���%��l���i��6�Iy�"�p!�W�b�J��Sܗ����ܶ6��݄f�i&��aõ��z_Hｰuzz'��k��6�9O�P�t��r%�Qd�|ƒAp����>�M���h��։B T�d�F���{|e�0f�$a��{�i)Rk��R�O�<wsYuC�IY�5P��34E�%X��#��9���^	�a
,s��b(�j%%�:��t���M�e���ݸ���qȕf�
�q�E�銘��~8���c#RcZ����QS1�YC�������W�8l҄gPxD����P2�6�+��voV)Wv�e��6a� �c���ܸ�b�]ƶ��U�þI,��>{{\ӟ�Ԯ¹��1)������oM�g��s�Jn�����^_mE���\L���D�G��s�wQz��8?:����`k��tu�8=!J�
��� b��3���KG��L	�8�z� �PK�t�lC>x�Ɛ�F^j������=�>d�z�B�S�0'�nm�2�+IU�a(�3�|��ͻ%֙�1qj�ƩW=Q�Zҋ%�A���:� p�]�;�v�}	�&��>���u��z��Ֆ{-���醦���Ax��U��_Ȅ\'�V��bu9�w	�Ab�u	�5�SzFT.�Ԅ~s5��l�O��o������,T%��$�Օķ���HA��;l�n����n�(hy3b��q��ﷻ�4���~G��2������ۑC��� �XR��	OC0�/nC$�I��^B��Bp���x1�JBe�So���Nqr 6��>!	O|�|�8����gN cy�<��D��J&�,B�D�iH9��3�%���G�61
'�e�T��
t[	S��D��=����8���N<f4���M�OFI5$mGx��{���R7�³k	�gϗ!W%��#��2C�0z�Zi�v�(y��z��/Wd%��@y��i°ȵ�ߔ��d�/:B0���e,$~�k��p�B�]����Q��Y�?����d����p h$���MSq�W�k�E�/`�;��TH쯂�N�����ǿ����S�Jp����+f=_����ݴ�Fzѝo�������:�)E��LN�&֌��{�n�1��M}����@��*1TƎ�,%���֍�]G?�|��1�p�z�9:��+J�b�Ӗ����G�Jv�f~�I����ټ$�v~ڿ,�"��mjs�����*_��N:��d�1�#?=|{�ڽu�9��e(��A�p����*�ۨ�����a�jv�Q;�.��7�B:�*h�mkO8�)�q��4�r�W����i8 @�	���\���{��yA��M˦�jDz�������1ʿq���=0�A�%%����BkU�����1�B@8z���@ԫQ?]MF��x���),x4�,+s��v�d}��G:�����@?�a/�~-W�OaW����s�����ϳ��$�:���o���h��9����g��&�Na����ho�� �ll�s���	�NO�p*mw�|Q|���`�� ���?z3+G5b�+6`W���y���
h>­N8>K�xJ�yQ`d��#<9�<��,��~��$/�f�b��Ts�P��^_�t�?��R�R�9�VB_�~?'G�(�s��X x��*�v�k�N�>$�[�pQ͚�D���ݪ�
�w�����܈	����품;��]h����N�2R��E^�������'�z�ffL�b��4�k��	�{}���G�rI���"O�lr��]�;��?8<;vߵ�
�Z{�og�˸G� Ѧ��V4���p�y�Ș��_���%����D��������{��2�5��{c=7��u��?9�F���J~8#�4TZ��z��)"x����_%!������aA�*��|"���
8"!��Jv�_�D��t��0���ņ�KК�1�֙z�A\�K�}�7�y��6����@Q�;T2�e��fM�	}7Y	U��UI���� *������BY��`,�L �ɇ&��i�}�e� ciu*!�\D�wԀP܀PT�6��1�'�5S!��x�,�gF"FiL���j<�|>��������N�q�-[^�&]&?R&�&R��N>ܐe܀�m�j~+�W��T�������+C�i3���;���>EقL�}K���p:��.
��K8g~���3�\=�����c��B}�$�5w3�9a���jOtc��p��P���
��s�p?�x�H��$t����k����TB�,��_2:��v�<נ�<��K�q3�見��2S�5H�����ʊzB�`M���v�F��z-�*����zl�u�=�HZM�Y�sc�����%�w]că�pb��D��s0D��`_�����{��W&X�y��n�
pdܑ�me���ٺ�R��Q󦉃��v�D2{xtq�u�L�I:�M�4�ޘ���A:�md=�s��s��Y�Y(nv*�<;��툚y�:T/U>ji����<�\��H>R`T3!��w�!�����d�Eb`dd��V���1f3����JJ������	���D6x����M�eVs''�b7�%��B]&铵$��6�ɓ���� :˺��V%=��)$8�5c��.:paϏ�6�K��:v�GgD��ms��;��|^����>õ^���6^����(�6�������=�������������j�g:�~ȊyDpkӃO�[�]�=X�r`�\��y["�m��zٞ�Y~�s�=�����-,AfTV��ʬx� ��V�5�����\�y~<�!$z)M$���w�hs?:J�h¶c��_LWߒk>�#���ri�<=/�:��OIM���T9O���׼�ZJa�NIH���o��r �}���xy�+�bEDDL�*ۣ�CC�cKɦB_�3�!��m�@6�n%��O*U��U^i)�e�������
�����w�.��HC�%�\�R��!�J]��XZjr*U��&���DK�k����^T'�ν��D.�k^�� �ũ����P�̭s����-��m'-�Eh��JE���B��㢊�G`��;gp������2H&0Pddd$O��\�`��g��[;=���a��]�X��B6f�ɕ�X9�,���B�e�R�]�.��������s�S}��h��#�C����འ�9�������n^^N�A��FT�k�?	���9|���Pbfw�p��4)x�����=��RP��(|Eظ�>%/kf����f,c��J�/����x�D�������l�#��2 ����=V����L�^����\�zNGG<�/�G<�xK9�ŏմ(�Ϣ��ClQ,���n���d.�`��ś�eai��Eް������s�3�=㯵b! �FU�Qn),@ӛ�\�sЍ�턌~�̑ܘ��SnC%���ŋ��j�v�:�`��$�U��-`hE`d<F}��X�y�hEc-hlą�8:9	ݼ��,=H%����z���|A�����!Q}�"A#$$��T{�l�a�jJj�F�`f�4i/$=��2�.P�Q!�e��E�z�No�Ҏ��Az@#Q��T��Ն��]`s+�8;-n�tum#$-^��m����>�ñ��.-�D�����	A}�HFs�!+�?P���K[�����򁶡���#s�1:X�����*���t�v��8[���!��3W����*^�k�V�h�:N�lw7u���oʎʞ5Y�ª;*��3E���- B���{�rmd���8����ZNl�t����;��Qҕ���d�B��$�b��!"� G���g�4~��2� �o�����\_qP_��[���^����HD0�U� P�1�>E����M�i�<�azT�����������Zo��:��;�!������e+	���[\��'[��R��ѱgg
���RRd�^�=�Dǔ۳S^��d��g̦�yV���������z�I*���8?F�)��c�Ϫ��� z�|߇���?�ump��8�r"!�p�ڊ&�Q!�wA]�{}�lm��:�6w���_Z�!��[>#��bʕ��c��Y��,.v[PQ �< | ����Bx��:_�Eb����S��B���l�jɭ���ҹE_����r3)�y�����]��N^�����ӈ��Ě�<%+��9���p>���������|��q��Mi,';щ������I^�'�^-'9"�	=JB�F�J#g(��d��Jr�mw�q~:�\��[�~u��Dӥ��y�0
R������Q�CsTf�^�(=+;��k^3�(�|5�S��,�^�Xx�};K�j�m]�mr���c5'�\m'A����P!����IE#��zv���=��[����$��������O.�^��Q$��J��^��	�_Z�>����U�)�(en̭��5��ڭE���4/9B���&X�˫�
qj9p���	xqo��At,���ˇ��:)=)��\:*�f�%9a��.֗<��rF��0��h_+J!;\��j!���1�t�����*!:A����!���h{z>���B���K쀱~2��c���wv���s���0^�%J��🜞^�_�u��U�hh���cH�~Wd���[I[Z�jؼ�������J��^��c��R~n\'$̯���!H�P��K]��C��'���Qo�ʁ�wfԬ�k����zRZ��9��_�?:"`�s���~�:GU �uѦ1�,_	H��j�,�����&��[��,�w:����aja��14�/��	�!���l_�^J��q�S�Ǐ���\E�#�F�-כT4ur��8�I��$W8�,�Ȟ��M��;ie��n&�6G��r��e/�/��:�t�T���Q5�5�P;4�sY��9��:��\��{|_s��~�5E��i�C%
�6vv�������R�T�MM��R\<<;p� Xؙ�ZYx�Ύ�ͨ��NB��n���&XBŝ��T*��ݢ�C��,U'��Tԅ�<�>��(t&����B�֢IJ8R4APY�� 6�����N���3�������"_M�-�v�1~�ų�B�{^5lҫUG���7}4�&e#�y�$�%�l�bC��A�I��6R�Oc�0Y1}�#�^�0��6����}>��|�   �YK+jaa!K�G9�i�����X��8O
?l������O����G=���|S����+�y�{��ḙ���T��O�[�kW�b7���<M������o��&��q tP����{4%`��s�W�"��Y��O�z�"�ݙB⿎γ]Z:c�o;�f]맏���!���޶���|�quh��z�[$x{�)��l�
ժ>]L�<��:x0����x����Ύ�[F_���,x�qp2�����Ip���W[~����[5�j�����J��YEv�a7���4%�R=n�F��s��/�#0�^9+[�ޔx����"TT[#�Wv��wGQ�E���K���k��ޱ�wV��.���c�z�~6b��΄体��Gk7��)(�Z!=���lͱU K.ujz:ddD������^�1�#<��-[E_LZN��'�D�n��:�_j	�!�Ǩ�w
����\-��ag����c��w�2��שIdX=��͐ֈ�N��x�T�q{[��u�V��mrPw�*Wj�6R���=F4m�7�q�W�G$�S�r#��Y�Ë��b�6������Ȃe�<>x���ł���'�j��e��ں�+�Z�0�͇H����36l�ʹP�K�����K�iψ�
L��'���ž��n+#�ϑ�%�_�t�3[�c]6~]�����|9�Z�	�+蹝�W�)�Ď��v��/����"���.���ໟ��L��p7IT����ʈ����%Ov��h9��x��p�K\�$8�É~(4��:aE�a�l\i����E���ՏO�;˫&��?1�� t��.f���@�vbUr�(��2)������k�1�c�������v>đj��J�y����]FfF��HxK���ܜ���t�:�P��w~�ӎ�T9F�n0�hUo�^N-I��i�x�b�D�`IO�3��) ^��Ak�x�d.�q5��nU�n�p�,'���H��{��Q���ߧ��1�I��Lnk'�\l,פ�0��q���7mH�|='��x~]�n��pt]A��\���3��m6����a2DvW�Y�dD��%���6����w���My_��6X؁�1����P�=����eh�O(	-�4�w"� p�|���.(��M�I9?r��"��EPG�@��I;�ů��� 87P���U�ڡ����=�c�6G�omaҾ^{]M��a��l+�¥�R-���[�$������nO;IC�7F�Z���]B����+���mwwww	��	�]�����ww�<@p��<�=|�����M�95̜3ջw����)������.�qs�I��\Ґ��w���"��h2�f��D�ӹ����=m.0�M��iæjQ�Y�G:)�q�FP�N3i{Y~S�6�z=�/�<�>_i��&2SA�{zu7�%�Z��]�05c��Wx������Q[˜�gFO.rp���r%lY���OG�ɏlg�{̗Ȱ�Q�}��I�0����|�+ɀ�_�̌�kt�"�Sh*�Bg�̣����2)*�F��L�  2�a�&�x���<�E��	����F
��z�Ϟ
O��<�J��9I�蚴l�@2��$�:���)4?tf�#s��rJ*nm�t_O�z�箿^]jhb�t��L�����~���u$�,�o���1���B������y�K��`u�������������s���jⲍ�����ݟ$eӅ*�Ë����-7|||1��6N��D���u��꺰�m=0��l��!�YOmS1�=��"�_r��p6��?�M�S37�������qހ��ɜKa)����Tbggګ2Ш�ÌW�X}�Abw��g"w�K���ۆ;d�E���o��x��e�M:%t��#�!����igm�����a��
�v���q�G��	r�|<[��lc�->I���C-55����8xF�+��?����Q#M��o��n�.v�5٣E}C8��U�T��8w�m��	2,:�[���}l~p�8z�P9��w(�yH;H`�DzTn���|�0����Bg��?Jb����e�˓X�y�`��85��_�p8l� w*��o�Ý�
'�}%]����I�f_L
� t�'��^J��s9��z�ږW����`�||�|�t�!�<�x���G�}z����Y����_?6'W��	�3z� ���%Y|� };,����Q��n�C߱k���Fc�*y����
ی�<7ڟ�����%>[�O�	��3�\�}�?o@�%$;��r3����>=�)[�}L��iZ�@�Sۆ"�#m�Rw�p���nIy����d�1w��
�t5�}�^��{�x������D@h�(f���;����%BNG���$P��h_�M��v~f�9j�y4�R���n�^�W����dK:|\�J��b)NZ��B�yM��v������2X��/�I,+_�i�n����E������6/��W�l�3����A[!��O)�v�h�s@��\a�>^�9/��(�e�H��u; ����|�5 Tq��E��B����
��J#��G
��z���ٟ�
��
�$O��F�-�*����MDjFw�Tm>�9���&>zƟH�0�w��$5��U�S%�C�� *���&��%�x�Vоb���T�X%W^�mj�k�cN����3W��2V�n�j�e����4�������(�Da�)��>�3�@A�s�^j�ұD��#�@���?���ٙ ���+��j.�L�/"��NcB���3���(b�:���.����Y-%̠rMmo�ꅂVߺ}ֆ�:�}��+��\5H:M�������=k�È���O�U�`��C��=� �Z�ky!��?	Ǩ?�[�����o>�;6겴�����:g�S���Q �� ��O����� ��ԸMm�/2����d�o�7�\��X�FI�.�b�Қ��5���&\�Cx������a��bC��L)��t�Z[I��|𶣕�\Ύ�P��iE>O]��!i�)��Ww��C��؉ �*F�h�?Z�]�ag'��m�V�#�3x�b��,E`歛<�(5���k@)�.�QqL�k_[��ɺ]�!>�)AV�X�k���r�HZEΎa$i|y�V�ى!�"Ob�V�>����mӣ
|�uj{A�Ϸ~"6���N-���m�c�G�����ⅹ9��B��r%z�D�����׏@y�K�(�;�5��Z����vϵ�`���r�AyU;~T!��`�ϑ\��!7���=�(Rk/T�%2�<lP}z�Ap�j��b�H����
��8��3��oM4�e̳�Ą�Uc��p�V������{�5����0�Nj��m9&.E�1��T��kyNk������'�z��#$�n��6�N����-�!F�󚠮iHV����e�,
���5un�y�L���cӝ����EJ�b����kZ<��w�"�˅��k�m]E�:�t�j���1ouF��A��r5MM8�?�$�LHX�5c"� ��M�&���X��Ҡ�|b��<��۟��fP�tx��S]���o���k}��Bh����'3�-������@+헝�e���M� �u%}������\���'c<���O.�x��!f���(�w�� u�}c��G27�IS��Uw��+��=t���A�,������	�W�����G�q�Ӌ�p�c�i0Q�O��]��о�T� ��md�\3���s����(�9m5��>IXd����Y���d�F����S.1o� $��|'�������w�Fi�H;�(��y�����%���������f���*��e&$���fވ�_�� x����Җ(��PNww��v]��s�\'777��,�zk) �	;��i�;�
��Ѡ�%N��J�}�v5�� �GRpxh���4���Y�H�]j����\vдXxt�h�Oe��Vs��q�?AN{k��iq�����+4nS��Y��ڶ�^��Rl�'�Dj
�8���?�X\I_>)����*}��K���}E�_;ֲݟ�N�|�u�w��v����i�Ae�n�,�_[�MY� ��*]���0����F�OvN�Xh͒"G�v#�z}�K����M}�x�:���:\�LޗF��g
��&�v��4ȣxq�p��s7���թ�����6��-�/^����o�d"H�}���0=/�ϊ�����[ ����o��?W$�/��O���qV�51�U��Cp[Gp�ى������A��=QB �غ��> B7����'�U�n=W����??�!�0)�ݸ5@�wY9!x�0l���1:H��l,�H��� �J�hn��~��������cn �O��M�4�3��5b��5�)2~,�	��`{�8��Jk"7��R:V;t�JW���B/�1?Km`Ѣ"�I���]��@R��g�S��۔����GE-�W�L4�z�%���z�����C$�Q��mthk�ed�[<�����4M:���H��7������(W�S������j��T%76J	:��"R��k3>}�e<u;�@C�eGG��3�;�ܖ��0����aa�Ez]A��ᛔܐ�r��%����TW�|
Re4�q���q@pl�e�͊Zs:ކ�u�!l� �N͎��FK�U�KIO�!���>�$R��gȺ�KL�tB��-+���^p-�&Rr��c����b
�[�X۶v?{���Ģ��,S��y�8)�u��	�v$�R�����<m�zs8QB��e�8�ę�p?hN���#!{�������&7%���zE,h�0�W��}�?�����.8��.�5h���3��C�C�ο�������z�ɩ"�k�f�2�!醾!=O���EШ�Q�Q���n?4�|�~գ����Y�r�C�~�]ÎF�{/�' ��.����-x��3���H1���}�_@��E���yqИ��+p�%��!ʏ�ի��}4��ݯ�W��>U ��)��v�o�z>c�U�W㑵��>]94�@��	�b�z���E���F��,��	�	�����I���T�8����`�?���/* �p�7B%�
D|t�&��In����ې��!r����{!!{�!x�4L�z��^�||��*�rz��E<ډ�7�Qz���.:
�<�ZZR"�����̃�O������ϳ�	絭nq֫?k՗>�c`<�M_K�^��'��vXwn_�d@�e筪��ϻ]���[m_ݞ���<�QH��9v�+�vW�����j�p�
@b߄|�A	��n�����f��2����@6����2)"ER�xe���;�j��s�|�Szs�C+��)��M���QZbk���(b&d�r��f�e|_������U4+x	�\X�W��X�"�.v�I��q٢����~�B./a�jp3M\���7�>�,4��teJ^�)��F~�7�5:)�4ut��D�#A��UU���F��!p�Yb����q-_�d^��
�	�p�T���sh?���`��tp1Po脚E���}�R6�SCL��1�J:Kt#O�~�[���E�ɠ�c5��2P����e������,�ාb߹�閭7sQ��!��Il�9b���A���*��GC$Ⲛ��� Bm���.H�P1RsZ0�b��o�J�@�)T{F��|��#��u�	ߣC��`�=�<��گ����6�򕶤D�^*�^y[|l��7>�͸���H���87�1�gd/����E�i�_6y����R�.��b���T�_Bp�4P�#Uf%$�r��aGbU�%!F�UoH�R����W�{K��8VX�VDL("Pn��ku�k�sǷ��Ya��m������BK|�Z���Y뱬(X���bnb�,�{Ǧ��ο�� �d�I)n°>�46�agt)��ށ�N�~�ƫr�Q/wJZ���}��W1�hѥ��EP�2kYfp�o�����^aQt�
<�U�	_�$%0�6�K��O|��Hγ��ư���n7X���I��Ƽ+�'	0�4~3��3K��j_�n2]�����e(��`"�s3�x��O��>�}���FU%�
¼�4�MT�e��䏇���q�9��*i���6����w�p�'3�Ψ1��N �P�g��lK}�F�����;  �K��	b��2���8D�c9��z�d<������?66v^{��U_�PbZ�v(^�*2e9#�h��Cgu=G�4:�x9�A�٧����ʋ�y�6�7Nz��B������q/
OF��>�B�%~�^��<�Y�=�|�~��E=9��r5.�@^Qu��{�Bmb�S{�/����O�&u��R�3s2�E���|k�sk\z޶g�Eav¤�����z[o��N�-�����Bo��y[f�N�L�/N�w�L�1}��;1l����r9�&u �Z������-�NN�C ��r�o�t�s��ح{�~`@�磫���:gKҿ�H�9۽=��i땧-��Ё��WZ?��j��9H�֬�������Y/M
�1>Np97a�^�IZ#�܂��)1��]߅\g<*�NF�i���ѥ���i���		��~2�D�)�|��O#�٥���g_p�!�{�?
xH�*mq���X	���ܯ��ٮ9$��f2vh<�B�x"o�&N�|����]H���Mτ"g�ھY��{t\�j��+݄���^۾{8lz�Ţ�����6���\ֈz��r`橰ߛ��a4���x3���w��f������|7��_x��Hm�Pj5LE�)3֣��bF��buQ���"��jI�t��a��jZ4$�_��L� �&��)@!��V���� jG���D��\W8�I�H�'O��J��P�k��Y��5&EJ5O}��XP>����4����GX�7�4�o3(=�<����&�ʽ��:�P�4/��`l�M�Ai����5��zϿB)�N�yWRKE�2��D���UA����!^�
��,�IL�U�L���AA�))>�:��O ͽj��������'EM��K��y\��z`i�]���jvB��I�H2���h)b���cU6�fI.:|���H�Qfǲ�ᗱ_P\`ɡ�q���J���%�#Ѻ��T�EZ38�����m���В�fu�4Y��;K��U�����<�A�V`5+�Z�Tq�g���-�0����|�3�%��sdddl�	�}��������2�H��� �/�DZ@�RH�_{j+84�vT'h�g�U�{�.��L���"|��O%b��R��x8$>�%��dUN���� _�y�4��i׉^����jk	K#���G���D����x�'����S�QP�G�zoTA>�S����W����Da�96>>�B�38c��J��P	
}��=9<
�P�E@΍�vƢ�w��	����D..[�T6��ZF��M�>Ԛ��30��/y���͸w����|�N�X�?��D���S�)���tݔT�t~�q�,P�_^M�d�q����p��Ɛ7�J�l�J�1�Fl΃���Q�Z�}sV��/��&���;�� ��V�C����A���֛LD�ԏZ^��`�v5�j�A��0��,���J=��>�I|^�]׿�49i #�yA��c�К�!���ԛ���mek29!��FWW��n-������d{�^C�
�M��d��d�L��C����]�[�3!@�������JPPP����D*����Y6�R�"�F-�O�p<�� ���ʽ�~������1��ߏ�@@A~��=�8��5��ɽH�w%�A���u�h�͝�s��8��Li+]گ��v\��Z:0���4t\9�e��y�;�!f"��n��Ҧ��M]co�΁�Qf�� IEe��^�%:���1���=v���P2�z���sR��,k�S���oi �7#�"5���yuS�����qk�h���l���b�2@Ĵ�/C=��͠�V�v%i�6�H�cه�Ͳ�� ��T|:I8��Ii�9�B^�ϲ W�����������#���1�s>����q�c���(�m�6��~����|�DlԈ��"��jw5f�ez/���;o�#K��ϊ�P��}<,''Ǆf��@�9���>8�6�儞�M�����9*﹗3�����������R��W��7�#���1���q`(�]��JB�_)�&�ƆtlJƒ�aLa�BC�\��$Zs#�s���9�ⵯ�3�Eޢq4Y�)�³6DTGe?`���p��ww+�����7Q�fЎ׻��1�9��%U%�1�ͰO����.$�Ќ�6n��~��37�9���t�w3�3�|���u�{��g���9�0����� ��i��>��i�D1DS�9n�!vc�:D|�gmm8���4�@�&Ad���dH��V���u�w�Avw�6���+	��*�Oϝv�ϞfV$�a�ӬT*;���w��3UD/0�Ư�
������-���a�������ׅ�i�O���g}B��G�DE�ϙ�t���u�)Ն���>���uKិ�	����ذ!�!���7�?M9��#����Ĭz��eк+���[��Zj�>f�\�9q>"�"|�`��UB��zOլ�#>�|�STDqh��������%��L
'ӛ�� /ݙQ`��������~?�*�Sd �]��KU�5�G���:�k�U�������?��!Z�a���Q��2/K�7����+(n��h!:�M��Ȱ�n����S:�_��Ϝ�'V������@����#�q��RQ���yО8�uC�NN�Di"O�K���O�:�q��ȟ��(����ơT���,����Դ�=]r�/(AHfFE<�����*3ȋ��t�<�la�;���XX��LL0x�������*���;!�}S�`v�@ Z v�U�q.����T?JL�]5|�d��c0,��PF��<#���� vX��w�\���=_�ؾ��ܒ5�ǳ;���v����"4��9@�	Qީ]��mJ_w��%�o�)�v���Dk� �DUB�	W����.ZY�0.������Ed����~ ����5Ʋ�e+�/V*�҅�>��2��Χ��v"u����8:x\����(@|u�����X��C:q����J;E�Ó�˱�]H��H�/��U�Ս<o�D���Y�t����t+��)Z{{;�W�do����ӞI2���7 ��כ���SnaM+h�wa{a��d+x`M�>M/��=`��|)�ʯ�1�%K����d�����g�b��ז
����]U�{PZ>?0-c|@.�M�%a\zVo���x�v��#��� �<�=�'�|�xUv����%�t)�[�Xֳ�~�'�I(����.h�64V+�XN�b̋zˈ�)���@!`��ŗA�x�:����`�;����贪���=�{���;vΒ�Z4�e���Lpp0drrr��<�N�{P ̎��zS�������Vq���PԿ�ݨ9B|���k��wg��3�TN�
z�-� ��7M[�+�����]��5f=60w�`�\6�B���K��y���	����w)%mIky���<j_ O��i�d�E��qU��@f��/��c��)����J����^$
���s��Zc����pq��Q��� �[�N�-|m
��x�$����<<vD_wE�nU�66��Ӕ($B��� #[)�뵬�VFCc��hZ��\��I�yV��>���b�Bs�ej����<9�P{|WP���B�͓�ǉq��9p9�5������\@O4��^�(�� <g k8�˧`�i���j'����)o?��(RM��f��$:����㛗��p�C�W]Ԯxk�G�n�����T���Zt�l���>�#]V_�hFae``>����kyz�{��v/���[��U��5���#�Ѣ�ȡwvv|�?](�����Ϳ���~gboo�ߛ�h���+_V^.�.b�����΋Ȅ)�0��|��X�~�p<-�Q���#پ�d�xr}E{P���H�ɱWH�6��Wi����'�$�Z�({#�/����!1�F���_���A�5��'>�!Htc'S�o�J8���H�)/���!�Tɸ	I���:�
z��ja��4����=};��aז�^~��V�ᗃ꒎�u�}���(L����Is4�D�&3\��%�����zZ���ӟ?�^�[���u��8�Pz�y<>2[4�8'd���c��`�a>]x{{{e��WG��!�9sF�}n�}ؕ1�Rh���BUW:"��X��A��d=�3k�� tLZ�${�8<�������F�E�)XhB&�'3�q��H�a�[�
M�k|y���54����z�������>�yv( %�؝cys���z�����C�����0N��sT��:���'��Y��*��GrYQ�_1��'Y���-h�R�����`���.j,$����I�U�lD/���M�!���L�'F��o��2B�u���T���j����5D�(ihH
HWNc��,�@�i=�tH�r'v�!�s�5�%�Y�f3Д���f��/>yj�&�8}���}��f���A�Ű�bئ蒨���K�sy�pB�3:���?�c�9]B�S ɝW6Dյ�:�G8��U�k��B#��>k`D������r't3x���c�������9��.�G~�Z͙����ɟ��^0��l��?B7\����/Y����s/�Ϋ���yd����:�.��10��Zn��ۓ8���F�3���|Dݟʍ�����S�u���p`;إzީV������	�Ԝ��w*�t��:*M�ƀ0�>��#�+��-@n�ED)�郵��v�9gU=ږD]y	�]Hl����g2�N��N,�QB���E��;�]��=���dȃ�,񙲑���Rj.PpF��5cr_N�����r|�����׶	�b�ֿ��٧��!/�^�Y��n���â>T�`pbbb�n>Eh����ˡ��(�O	�i�='�?Q`��D�2��ǑE��ڧT'7Pҫ&�h@�/0�PZk�<)�ӎ#7Ð��s�b�(���&"���� �6��'3�~_���U�,��h�f�!����8o��`!墁Y��H���X�Gd3o�eA�Tpq\���f=�j"�j	���4B�����{8nr1�4�.�����#��V<��s�9]����O_w�v�](�S�[���\����P�x��f��w�VW ���� Vw��}�^a����DJRF�n�*�0Bz'p���s��}�{#���)W���S���>p(�����;�k�%�<���q�œ�kz�!�^�8j��6L��*�����Q�W힮��<�R忷�K�Ka���^>����G4��lAϝ��FC�S�� MDFA�sh ��?�ぁc�l�����]g�$�����'���M���\�:� �1��������$��O/º׺�[H�]U��q�5�W��V�؋�,�tO9ִ�c28��m~2Q�"hHl���D��r��	/��Ps�[6E�c�����f�~��@�5i�u~{�7;���s�o�w�A���v�Ǎ��3n���Y7�>��MM�fQbCet���K�1EB ;��([}ٞQ��<��턉���)))��J�0�<۽��3�I~~yYs�.2��*f��_m);t�etl;D뉮�U�r�^�ȺsV׃�I�M{�`��0�k�t��ž7�'@�߯�ds�y�T$FR��*J¿�L$����E��%�B�N�1��_��?���=9������R�ԑ|�b������ѐ�D5��M��nGjU������������u��T1[B�eڟz�LDQ�ז��z��]ҡ�1�Ϋ�x�tʞ��_�����ڙ��]�v	�V�P|)N�H��<��p��#q|�d��2����t�gl}f*�j��X��������gE�%��Feuu�a�0q��W �aX��Qs�>c�f��p��:(7��-�w��59����JIO�a�"��^B����y55�>| ����S�?�ճ�V��Ċ�z�\��/�b�T?!�rN^E�H�Տ�a:I� �i�40�@~�Xŕ�d���Q�hs$�vb��Řl�e����)�w�y�Vg����K+�HZZ�K��j���3�X�SѨ���1��j<�(�u��2��� `������<����4�#FM��)h�T�x�g<�����!���)�F��!��z��Ly��QU%+M���,py�o��,3mS8��I��JU�?=�4	�8��"zLZB��W�:x�������q����^����i������)G����g�I�55!A�5�8�%S�+*T4���p�u
��-�UPPf�b��E�:<��(��jf�$�/���a��&�Kq3�����^��Z���6������� �u3�7���"����$lmTg{�OG���e��Z�y2�y�_��Q�q�qwx��$JB����n�+8�xՍb)�}�gT�F��k�>:w����Z���������w��ON�>�!�k����%�A4�=�����Ynn���~"df����(�#���؍Fa$o&V�3�	F�َ[��9���!:
��yo��y��0���|g�3���u�*�N�a��>Ƽ9/k����sS������3�ǁ�F���Q<h�.�=�nOX����y���;�'�{�	�u�]D�K�\$
�e�K��Z�*�z��j7! 5l�n2��ď��^;>�i���21_� �j�^ ��VS:7A^��r�3�7%�?}[�F8\Yʺ�TK��;f����a���%��5X�C)��{��_p���)�HG`��S�ۖ3�sE��[�䷴I��������Xtn���"�s<�҆��(��|=Q�!X�ń��q�l�����5C��tn�b,ŞE�=:�]��:2e�Qlh$�'?~^�-O�CeK}E9l�z2�~<�j�z#�jopF4fcbddd�^�J�_@>>���=*?Ñ��tzG�ab`�:;C�
$�2Q��4B??�o3��`�����4��E/8Y;ڠx~Qp�~{�#][�s��-v �Ƙ0F&��6;&k�b`L# �||�F���U�t#Q����ǧw��:{�y���-KjXtʂm�liv|�c�P��&��Ev��	��&N�ay�o8��*n`��.��#5ޠHxpn�I{���`L�Cx�����8��@�/v�Ah<��i
F��\�|,`��S~:l�T��%Pr�*&�:P�2����ôQ���j����[R�	$%���$͓+Nc\I_n��me���xC"��w��)����,���h�Ca����QW���8bU0jfY?�!:D��������=������9E:ં�H=5U�R3�>�����`�ʼ�N=�dO(ñ	��q �RkW9.�4]������r�����f�����e@W՚հ�i&�nEݣ����{��ڌ�2읙��������^v�)�9��n��y�h��Q_�-(��fT�5�Iho#0��x�'�n�إʦD��L�:�Xr��GHt��c�U����Z>V�~�ན�<�]E�K�r��pi����
e$�4đ^��K���js���>*�Wڕ�B���w�
��I8o��)0*���1�t�eX��2�$���/4�t)�K�_q߃5sJ>���.���������jXW�?�>�D�ؠ3t�(�"��uC,!r맰��
���UH��,F�g��\�R �Bk?}�ܓ����|�N�������_��T��o�5ۢ�(5�'"�t��U�[if�^B-|O��~�?�ǊzW��AtX�j��:��:��-������8��׵" j�(���Y?��鯇�,H�g��� -�����˞�j��Q�^M������P9����:��3��vG��
��*��r�ݦ�z�D��;V�.�ipl�R�zD��΅�7�tD�w!GH,p�eT��/v@}ϸ�O�nk�L�&��?�k�S?7�}<Ԩ�Y�XdN����l��-:�����<̾�"��G��%t�;r�̇�fp�V�oK*�b�;.�7��Rih�Ǧy*����_j-�U�@,��H5K4h�3&�!V����P�ˀ��^��"C�Jo6xć����y��Ҿ�~2mr��s�^��r?0OR�-�ܤ��;��9b���Ft�$�\��F��@L���J�M�JC?A��q/�7�7���6�ժ˥j�ء������*����M���	��_9-�P���-/j��v��Ư�����Z���<s�kD(�@��p�:}�5�sE5���\"z�V�B��éu~�Y1dTIj���Nv�v}�f�</�nO'8H��.�g�}�S�6_�L�Q�I���c��O��;��=�:k��Hd���x�yu7��;LKe���@�TӍ�۲2�`�4AZ����~�,�;=��Ǹ�����%�	�x:BZ[�.�Yp�Y�#c'[�L�/AJ��H�g!%{�޴���x���	�ZF��������ŧ�2~	|ݗ;�Wq���'����&���)�=��&숃˺���r�������kד�����N�;�<�]&]��kؕ�������j0Mf�Ө����o�+��_7"�6ɪ��>PxN)����z���=�W�r��<�:�:�N,-��l�V����.a����ŇCR֭]�Z�v+�2P<�SGYƕT�����d	�#�;<s��nu��/��(i,TA��P_	��y�jV�`9(�9w�|nC��7�깂:<�y�����F_zot����(�s�a�4iJ9�{�C���fe����G���;��W �=s��o��pD��{q7��oGz��>\Xv�zY���i6#��6�}M��7C=�X�z�i�}	�L��C�,�.R�@��I�"~Ґٰ�s��mU����:zh�������Y�Ы�Ԟa��fD��$��r����}�*�~SQ�Ϊ#� ����9�(w��GU�F�L���9��'N�f������߽�����[�ڝ5�CPX;`N5�b�㢻u�ek� �*��;��%�����j+��z�k  �����/M�a6���U84.��g��/�{=�	|�6yF#w��2z\�ş~�T��R'��I���Pz"�AH$�1�H��/�8,ںF( �����E�O�)�^�6�U�	�;��k(_�M�3$J|e���d�[NVd�-|]k����u5Q����s�)���P��;uD��Uj��5��v?���n����ا��[�RS�7|A	��1k{Cd�ޓD���s*4L|خ��q�؍2�cC�V�y:��6��+����k>�b�G��)�hh$(��WC/�����Y{�,���)ښ�q��t@Xkf:�i�P]{��o{�*:�|@�?��>��:h�*�v��l�h����cGZ��տ 3�'�,���F�Q�ۼ�����x^�p���nE�8���c�`m���Y������X��C{�ř����[�&��T�����틳X#�O"��%3��+*X�㵩�ڿoۏ~����5b�`D�U�������<:���[�x�^�{R��.�����ѹ; p�o��5�����WO�����Yv1f�_��,Hx���V�f��������x�tL���2-lX>x�W\�^�M$\1���>&��J�L_l��&�f�'1$������=�P��0��~)]a$.c}(����ȻmV.o������v��#J�!����:��M�o�o���||	f5n�B7%����i��}Y������iv�MD�7�O�V,�Q�4��mڢ���@6��wֈ$D��&Sjm���1������`9�S��l���1�g�'���4�$� ���wK�y[C�~�o�`[دܱ�~�?��D��y���j*vԜ�e�t��8'��s���J5~��޲=v\���~uI�K֊�O]@����u���G��$;�x���_�!Z{B|�������TPK�$����΃�y��d�i�:��R�O�xlwzL��S���~b8��]5���2P5��b|���Y��lX�ST_K>A�Ɂ�+�
]��f�
��FdK`u��|
f��hg�B����l���E^_7�[�\��xz�H���:���^j4��k���s�g~f`N��Z�^���´��r�G��JU뾢��D:S��;{�4�]�B� �3���p�[Y��&�j۔Q����O�VyT�yt�e�x�x�jl�3F��{������ߥ�s5ǟs��	���P{�ޢE�c��9Mf��z����f���/�[+p��A��Szaw?��A�pa���n�ƶ>���i�V\����o'�k�E�W�&��e����)N(�d�Q�rL�Gk_5s�iI�=}�載`�`�E,�N�%��]tw��矶��Z��_&8���<g��[^@5�I���O~�t�6O��찶�\��=}���7����uq��o߷t�B5�z% 8?_Rk�}��)�c�ZG�1�����`=̇G�\�=6-����"�?���[��ݗ�h'�/�M�_B�h�N_�����A���Uu�T����"
y[Ջv�iI�w�b��g�堙���g>Oo��kM>ʇ(t�����t9^�"�k�52�o�y��?`
�?�q��K�)��S������.&<��0]�KB��L�Q�ve�Y�����ԸC(5�g��Y-fTpN�@79������xg؉��%V������6�=���h)XǢ�=��*P�}�ir}�$b� ��e�\�3a�ץoG�/�R���/�'=����9��ɓ1l��N�X���7SO]��j�p�6�j%����2�T��W�?��G����I������bF�nzH�';�!Lh�i��:m{�D��M�,my=!*y��x"�v�/�:T���,�;����4���YҞ���p6�mo���o�z��[+��˱�&n^����M;���/$0��B�b�C'[}�.��Q�2���πS��j#oB8���N��~�S�p��xǒ"K�p�M����XjD�����6̑[{�Q,����M�����<3�\���@|����������N��*\�(������R��gC(�J�3�d9�T�~�U2�l��/D�?�5w �GS��{x���69��۲Vdol��d�qS��P��RCX����HW�o8�7�=*	����W�>���b$*wpr�}_u���QE2-�Y�z*f���8V�Q�&�f?���OǗ���d��4�Dsz�%Ζ}�Af�_/�#�S����R=���+���F&��1fx�YДe��tF�FĂ�/����:�ܤ�@=υh�FF��=μ��6O�r��}�Z<D8�S���5'Th�3-��	�tǾ@�d����LpWD��ՙ	��)k�H1�	m{��cWr�u_{���N<��+6�l��xw�[g%Y�k.�VR��V��&|�<d�Ώ�U������D-*1�<�,#�7�t4�y0�a���ʲN|u�lI5��lL��~����ͭO]	���S��>��V��=E��m�Z��}68Ǭ6L�}�����a-_$F�3��W�Z�g� ����+-�T�$R&xH~_�$�@h�!iQ�e�Z6v3GJ'좊���WҢ��m���{����-ܠ����{�*��Yˮ�:�)����Ӊ�?��K���芡��ۭ�,����� zy.�@� ��Gs�+C�b����[�hf�x=qZ��^]�'�/�$����}Z�_b=
�I�ژ,}{>`���TT�cnКɃʿ�|n������L�R'�P{��o�]_+Z�AQ��7�ny��s���t�Ã;���!�wwwww����݃�&�������'�+����a�T�޽W����>5��b7���Z?g�켯>m}�$;l��G��qo�O4;�E#>��r[>��w_�h��b"�Q�C [��[ٻQ�D��⯖W%��u�n�h��	�O���G���D�Y��R{ �,~p��۲���z�Ğ�W,]��=w}����{�f�W�]Ix��6���U[��5���gN�!6=���D���\��� ��O�I�@ű6y #��n������60P>�wt�F	�!�j裂(�P��;�D���ި�������\Kџn��,��u.]�q�f=���=7�fQ8@D��A#������t�}rq�U"�	��1�/��a7����l'�3�_�ZGn{y؟?H�}o���u���@�/B$<�r�m$��½���Ih%ڳq����%�ɢK�43�m�y ��+����m�v�/��X�Kc LS�=���hIG>Ǹ �j���>�Vs�����-[�SJ}4f���w��ݬ�00�&����ȑcH8}���B���&M�����&D�9q� �~�Ȣo*j�Y��df׷�K������zv�:��]יh��!�z%���)��v������p4��<.��YD@E�(}j��y�ג3��s� ��d0]�q��BF�tq�XSe�s���1a��J~c�'�]l}�=�jh�(�n��j� ��c ����$���,Z> r�Y����m�?�l��3���$ad�;�aQ�w *�e�>��Z�� ��~R���1|dr�}�)onx�?��^��Ȼ�T}߽��+]���'Տ۱�b��s����!���m��(���pZ�u�e�H�9�W[�F�P�������JB���N�3����7"�I��6Cn4y��n�G�8�|�y��|q�a�.�y˸'^��Ԏ��{��о�VB�M�hb�`��}2�6SU�u�1 l4��h��%�{�>���2m�Hc�l��F����F9+���̲����d 	~�̫�3�"ȝ08/�Z	���ʱ��W�OZ!.W������W�Y��I�f���H���@A��T��#iz�k�t$�����eVPh�y��\ �%l��h$����?V����	�j�B%4���z>�U2�M��9��XI��i��m\�x�:����Ā0��m�hv����⺦��O� �]&��~=Y��f7��X,�:s(��&�i���؜��#��:��"�*ǫ�OK�>�O�͸����ZI���>J�݂@5�x�6��J�^J�\�K"�1�e�M�
c0_�j3�^����V_�D�	S�7J�1R��ń�]&D�q��ڥ��jrw,��t��|�r�������sPҎ,(�u&�	�c�DM�j{Q`���wt��a]i����j��[Eؕ��+QVÎ�Lr$U�~Qm$΁�V��U %"3#��o��Q$.�Ly��bƠ$@��2��l(!��a���;�c;fN���}��'��LN�ciwÁ�������@G��~�jO�7ƚʬ��P�>.�_�r�j؈yz5,�͟Vw����$�{�T����Yߖ���,#"�l��m��2��o!.�ӌ��G��,rOW�2+�P���jԦ#�V:��j�zЮ�R��}��&�(k���k���\�s����5��'_i��Y7�mI�R\/9�F��>V���>�P̿����x5��	0�	(�{w�$	��Go=��*O�y��>j$	`9�"M��̼p��D�ˋ Q�Or��QR&���3�â~�p�d�V� 0:�Bo�[�h
>4{$@'�F����|:�>:V8K��{n�׆:g>qz�By`�>�^a٧+�q]����[�G�GM�IR}��G]8Tl�����ߤh(�Q���U�"a�1�F���PB�p�e:+q�j؅J�����Ћ++G�
Nf�Y�5*�3<&��p_tɍ���U�*��mMvS��k�>��I��u}p�
n�Vt���Aa���]&Lц�GC�:%d�Y��;��˷�������{w�z�
��O\ywJ�o��3f�������#���#���pj�Kt>��f��\�P�X�L���zҥj���YY��1�,��L�4f�cG�͞��!�7#�m���& �`?)�!ڜ�1?v[�,�Y�Z�
�<�ƴ�y�:t�7��/8k���M���p���**(��CF/�q}���O�)ID�M/���Ǜs��A�&���Jo#$�]��($	��ݻY9��$���n դ�IE�sC�O��q��q糶�49������� ���9�?0���x���������z�N� C�Y�p�����I��~{wYY���r̰qд�-�K���F�ۥ����ok�߸�n���ͬE��k� b܇�%!��OIR�ifb�]� M��F��c�
�T�fs�$@�iXM��7T<>Hy�2�d"B�.T�~���;�:[:�������3��$���H�Vpp�]H���=%wOFR 0ٰ�
�u�yv7��j�#J��Ng��I�st�륈De��ԝ�L��X$5���������� 9 \�X�
�Y��0���})�++D��/l��֪&̡L�Ύ����7� �cD	;m�ޖ	w]��)��%׍b׹ݣׇk��
�\��e�� �@�Rw#33Jq��Y6vv��Y.;Εxq
J�Z@A�p>�|��g��"C
���#@�<<��-2@�k��y��{�NdEx������=2[��>�"���U���\�;g=��^9p�.Vn^v|��U�*��v̅��SU�)E�$.j��g,Dl_�|������(Oxb?fL/�s.�����jI��=�����S����9v��1�~C I��uWǷ�g�ӎxZ�����fe %�����`Aj�s@��8���&��#�ƪ�pnC���tQۀ@b@�'hȓz����_�Rc�����\��6��~�C��6�7jY����\�0Km��^���o�FG�'@`��~E>2�U������n����?�;�f%,l���OU����_����T��~2����'�AG���Kf+ʣ�ҋ܆�cS�����I��%����j�f���������1]4d�N��+q
����&n0�ҙϹ|sӃ�̹�tQ��V��W��>6\���zCy7?2�rn V��?B�ў���aь��E&͗q��]ӫ:�@��5?	�I�L���>r���\se����q����@E(�`Xf�J" yQ��j $u�}_�t����QϏ���ŝ*}X�H��e������&z�eii|2ev+`zj�ב6���j�+�έ��vB�iw�&��s�ᣀ�H����'�q��Y�A��}�YXu�Q�v�;A�x�Y�����1�f�+\ ���	;,ܞ#��+�˶�}����6�
1�t��Z����M%�d�ڷ1:���2�2�X�W�#k �UO�rjk�*.�fJO�
Ñ7W"� ]�0�k-�= P�?� � �O�=��O���cwY��6��̗���R��V�Kx�h�[=5�Ѽ ���>�d_�+�Y����Mӄ~sC����<�:MیnÅ�$��';U�����y#6$]t�8��4kP�R-j��g����PWCS�����;�����l�<V��vsJ���b�G�)��h
?����MU�)r��P~92(7��xbOԓ�7���(0��2H�|$�Җ�i~�����^!e����	566����O�~fH)P��O������V��6�����@�f����Q]�ME�ܑ��η��L�A�<�Rp�Rm�Q�@�
LQW=I�T��|��y�n�����yk)v�i.&�s 󱷋���:�������tA3��8�>!*�Ĩf��p[�J��N�Ξ�͞6���t�3e��#ƚ�T�I��m�ًf�v~��C���w=���Ҧ��ug�C-)݄Hv?SN:_�-�s�Ud����~O��ܞPp��z]�(v��Ŗ��ǳ�s*��<��5����4iVm�5���'�����C@t�JA�Ƿ�-����NK�7׭���Y���eS,�@����}��$3@�p�_Y�>����5�����5ɢ)L��\�d��3ڣ��� ��ᷴ;���0 r���,te�N�8�}?���5�0�5�2��} �=J��y=�y�b��vM놻ǡ*e��#����M���J�40�	�9�4�žzt�A(��!���={t'�qfw��{��M�
�-��_m#D<?�1��MpTE��44�~�`�R^p��I�w�\dB~ȝ=�Wý^���c���!��+�VQ&���bv�1�����#b�,^����t?�ǆ�&�a���K�WE&&h�l5����U  ���q 9U_�M�`
�ؚӑ��'�]L�'aU��f��\�����*�'�2\`^`$�w��>:E4u:��-�L$�F�--S�6���z��~���!�A��=����)xʴn�ɕz�����0P��I��~��˥\�n�K�4���`� ��k��e"z���{���'��͆zW�A�]�N��U%�O�2�Z�Q��(b8���In17{�1�G���_ T�yB�8o�L��s�g�!m�B�����Hq�E�T�_Ru��t{!o^����ե�G)Ä����BA]+A�Ct�M2pE#FX����(~�˴���s�bQ�-���׀� �
�����?280[;�c�G������
�h(��p��D�o��2���U��T���T��)�e�P��\iݹ�S�`����QN�"�Ӕ� y�ڇq��җ��ZDT� �'���őۏ'��� �'�L��^XȄ��cFQJ���5s����R=����	-��~@]56��.���bd&��(fE���Y�@��F�@ ���UƯ�#�.j@��
&4���w�߽c;��˓��'-c�w�a`BDb,:a�?�3���y�W������+�*�'EJA�6dEQVW�a�Y�(�aN��j��*�~d2�t�h�R*ּFV�W~q~�HOvx�I7��'v��i�0I��`�U��A��7ɿKY ��q��~'2E ���;�EM{3��������&{�.sƮ�e(��@xT��@�C������;��4���SI%WP���F]zZ�5L�_k+z��N%~�3A��[�8�{M܂�x�k �¯2RpJ���X}���XW�d���e|+�W�����_w�I���/�=B����˩�C�\�*���ږ���by3�œz 1l�@�4�@%2Z�a{�|�gU�}]�ݷ��$D�2DD�;,�D&E%�^m��wD:��u��m�����&U� �'K7�����23�z}5�h�(���^)]��[��'`����{����m����9a�j�՞�����/���/��u��-ϖ�lQ`��|���8��9�x��BL�P�4�.�x� ކQF�JN�5�U�<%죙U����]�"�� iN��C�5�n�u,ځ����.eD�˩���y�F[����OV���TM˄ԎO��]�7{k��T������Z��I�4{�!]�7�k[s�M��0Nd��/|>�k�G��1Fs�Q{�&\	'�
����T���&�_����:y���:�9���n[��t���5J��a��dS�XǼzA��{��Q���!!_��?����U/�����!���ҵ�U��Ϯ�LmQ�ĝ港�/�T�ZoX3�h���M�
�(��V5g*�iw+��Ř$G����P��F���`t>�`��;����A�奄�����t�x5</Κ��KX�z���F;|9+���*���f��	k�e��W�2�Y�ʺ>�Q��x��.+ף�)
D���Sz�����fP]�=O���ּ�;��1-�;^/t����W��<�w�=`"J�4��r������!BMA��B���������J�$w�	�?�iW|��a�kj�x�j�EX����9>�������7�i^G3��i]�0Epeg�q��V���p���փ��%/�:[eg�<��;�o�7�1�E����_e1n/��5S�V���*1���ԛJϹSB_<喚2�S�"��>�!؂8�9U:Ci(~DEZ��V���k����W�,q�R$��u����62t?����Y,�����]ɐ�e��u1UW0�m4�QR��������k満�/R���	�}H�H�������߀�i��Q�d�0��F�"
�L��a'b1 ߸�|�C�I76Ҳ��N\\շh 0����qft��O�~�VOar��Qj((xtt�Y�=���H�Ï(���0Y�D##�9?:��!�w��������kr�Y��
�������HD����u���p������~XcM��ˆ�]Ƣ��5��k����v"��5uT{��Q��_4č��:CŁ�I^\3��b�UA\�W���0f_M>y�_�c���?�~�byRc���Z���_�m0 ��c�hR�~f-w_[���m�βC ���f����w��z����Dx�4��9�¾j�,�h���a��`���pH(��"8i��A"ZW�*��&7��|��Q�D����L�23o�D��M��D=�xFˎ`��N��Hw��8��<�B*�olɔ�PT�l��Zs/�0�-�-�}�+6�-17�ˁ� O5	H1��B޸�!Vm�+�]B_Íᱟ[����o�Y�5��o<@�X��}@s?r�ˢZ[3L�#y�hzV6��.�`�c�NY�#)Vp?y�豂΍L�K��8%:��S�\H�l^IЖ�(��Iu�6�f����5�`d�JY=��P?-��Y�ym\��R���+\�O|����x�x���"����p������o3la"P�����/TQƽHIΣd�W�ح�Ș�1U���Cd�e��� ���`�.x�B�U_�b�9��Z{����y��z�z�.�d����Y��@�?G
���u|�VO�CUGЦ$�*Y���}{m�����[�ǂ�;�5$Hm��ڢ d�}�>D1�,`6���3� ��(? ,�h�hvˢ���F�e]�aH�\�������|�,���
maaS��<y�IU.��������0v5_���ݧ�d	q�9v$R|drqӒ�x:A�� Y���1��(u�R���.S�:��Ҿ���4W�Y���Cl�EVF
�U��^�,;�a�����"e���~r�D�X�E�0x��1Fb��xvA�	�֭�&�R�Cʫ�I��ԏ��C���h(J�<4?�O���,�t�90	�,�3n�SVY	�f�����v� ��͏+)��DB��:�0x�s����хQ1t+�V�YVl.�4fO������RQe/�w@��2��@�ؠg���s�s��|Q��y�PɊ�w^9:�ve��´�2z��2����y�߁���9l�0�K؞��
˜�,���ۈRW6���:R!Rd�qqj��IX1x�ߧL��PN8#o��AV3����4#+}��`�iW������ks��z��L�f��PR�A�6���a��zl�1iۡ�[9NଔQ�?�
6�0cL���y+��I�jd<=xTgt�	�XS)�����nI�Ľͻ���(�P�X��DF&�?���b&A\=���S����}��4��s6ZA@Cq�����S��~�ȧ����}�y匑�"K���䁫�P�Y+�%y��gsU�,y��'W���	^���+]�A�s+�(;@h[��5�]��-����[.����
����t5��a(CL�^'��	kL-�u��$h��#��j��g���:{�p��h��?�ׅ��P����kIL#M1�Ч���g��[MG�f�:���3�����]���6�<��E2
v�R@�;�N�4��~�WM9��PK�qG$�u���0@�`3Y.%7����zt�yd���-'n����4bO��A�Gԝ���*pG]�tD�a
P8:�@����ɤ�mg��@)U��	�^�ՉJ.җb3ԟp���5����[q�6G.�6�&����ܔ���Mn��������M�dV�y/�E�b�/t9�$W��Fz� �+�=�I��v����H/����94�TC�}���i������{��G���6�{`�|��W�	헠����!/"i�c�>�*Z*�w�%Vk�
q���d�L��{p�n��`Q�C���4��dɠ�Q#�{�s]0YA�7�)!na���«>r��bG�KX�.E�~�1�+ �O����͟j��=&�j�9W��D�|7��Ф(�����s/t�
NA�9�S���)��>�[�lu��o���ڍ�bo�wV�?o�/�{�U�����z�.��>̮{���5E��n���"7Ҧ��r�#�#Kj���韖���P��u�˥�H�v/_���uh����m���t�`hP)�#�]4�z����{<�����8���V�}�����p��4��c)5���HfQ+r(!�J��</��O��?��_��;��
퐌��w��J����i��.��H�X.z�<���U͆���y�����6	��m�K��.��NGc�%=��u������ �t�%7A��ZÍ{6�Q
z6N�`����@�J �E}�L���jӛ���,�㬛if�I�T��Z]tb���v���×��ڶM��9����=��{2$�����
)��|L	�_x�8�ѷ[9k���Ev�M2�h
��-�5����Z��KpyE���t��C�c]��}��� �A��/�>\�����C*S�ʯ����)�;p�~m�A8u桝�6£��W�Ȳ������T�t);z�,+��O���������SC���iנ��JE�l�Q��9޶8��{�wͯ~]tf[�e���f	1�^�)�z��'�Vm�
=@^��g�P��6���^��c�:v���kt�~$7�(yE!�$�4& ������K��(����ӳ1wo�C�}�j�'����!F��6s'/���FًJ����_��	��#���7�E| p���kpr�ә�!<��I�������8��R�v�b/��N��p��	g��9ݔ��BW��B�-��jQUɡ^K���ij��#��ֳ�掠�i�P'��?MmE�ɬz.H���{
&M!V�Ԁ�
�ޤJ1�Ox��y]윪��o܃*�q~hu���G���h�_��s2��I(G�~]p���l95g�ѷ~�f�Ao���d�}�����t��Ty�d=i'��
D�����~�Ot���m�5�3C�0~�Ӡ	����E_��q���������J(@X���C��Q��������э�RL�{�pR�?�m����z�	F�l�<g��Y�:b��z�,��z��ϟIٻ����W�l
RfC'N��n��l�O�|q=���9�'�_(���x�E�^��=�}����)M�&�>��V����pc�}$����]�,k�O�f	��PHEz^��k�%|*����	ȗ>=:��4y��9m3$��+P�tH��0��F73ڕvB��r�nZ�Z�?A�R�۞��~-ׇ�����hQ���/D���F������c �4����A���a��*"m����,���r��3~K��t��IZ�.�^�5�d�r�y�U<�cx�-!�����³���/��ll���[�;ރ+�����/���h������/��+S��u��8���|��vNS�����e�K\	^��]Dq+�m�A-�3�1�8��H�hd�����'�cRIW��w��&�������Kb?�^M�5mO_�?Ś��'������I۪�������<��惋�J�
����^�J�q�[�Ŵr��B��[al�r��Wv���ۧ(sי)��?~��M�#�U��ik�*W��_^+U� b�F�#`�n�s,Oy�ӽ�����r�K�"ZAʼ��9(z��� �!}TQһ�K��n��E��e�@�y:W�������~��{v����n�����Xyϻ�3�� f�.�um'��ٿw�����7���Q���UZ��߰�������b���c�#qt�
�~�&�u�&�4b%���u}ǣ��:��s4���Q���ٮ� �1y�+�s���[�<��Y�Y)�Zc����*�᠙��� �:z��N�;��Ңc��ID��Ƿ��7Iy܎h�7�~�7GT�B�q��D����z|)��<_��O~{|٘�!e޽��KB��9�*�_�'���.�|�d�NԺe��0Ns51���S׹���ϫar��
�T��h
��h�l�i���y��4q�8w
^6��o+#����w����V}Z�	k���v���Z4m#���+=e�������̪#�#���/��|}ص�4�x<�G��
T$|f�s�z�2M	���t�����%�����Qҧ�A���MQmJ֣E~jаF,�;��nq?H��K�f��#k���.��E�G�p��ǿS̢�}��4�=�%��9�'�sEm7&�n�MP)���M�nF��p )/�(~h�k��*����FP�-h��B^D�!��ɧ�k���� e���l�A٩�7B���a�N��_�Ub�f��l� ��Oo�\��v>*��h��.��>?"�܄�b��y[�p�����Q|�(_��7����3�=�?�iy��zo`�i�Ik��:1��h���Db��G���8�_��nΐ%���q���������p����:� S����L�ó��$�?����hkϻ�x�󬭷KG /���U�M�L��q�8j��EHv������k%��X�>N��@[L�fRB�J�K"8��qM�*Mx�����mܫ1i�a#�i���[T҃��;z�o��j!)K���1��f��;���U��t�>	�Ed!�i�U�����VR���aV�$2�@8��+}#]u�-]n�����Y��!O�G�)o�����v���p���&o��[�a?ҭ�q�1����9���N�5ѵ��C��6�Y>`��~-�[Qn En�O�[&��I�!���*���&f��?k";��Os�Wr�x�/���DL��7uC�!�2�yLa���pNU���E0ϛ��T�޿�*��>��-x�`\�}������qN�x��	,��ߧ=	�L�E��u�p��-^t�Mw��f����ز�]���_G����"�E�C�Δ��7Oã��+�J��?�[�K�Y�4���xp��ٗ��[a���R#��xB�/R����I�/���L�Oa���&~ ��j Y��C_�HH��N����2b�$�oV �*3��s`�Ê�C�UW�7,�x�=��!���?���jzlx��L*ZK
�+��bv.GZ�-F��Qg�e	�oƧ+��+[b#�(�C}H���6K�)*'�gb4���CA��q�\%Pj��TE�ol�����D��(�����h������i��� �m����14QV��Ens�����à�v|ﮠ�����G1�����+�������}u5��K���ٛ��n�����&�ؓ�odu�&��2�H��%��� �!�p�.:kѰ�ܨY%�u{�3��̰e1Itl��3��k?��MTa0���. Z�n����U���p�T�=����W
Z>
�	�#�o����;-8��=��&D�(O����V�� ���ϡ��E�I$��1���CEIt�z� a�r���H�F��5br��.����Q?���
�Ec��:�<�"R�zC5Um�p�Cd-��o
��7;��k9~����6�����փ�]��r�C�`\ �'����`t%ߟXV�kUU'^-u�ΝOi�n��Yx����\DT
�dn�U�,�X��]s�FN��$��!`�;�q-➛s����_�w���mMF��տ~R�ߠ �ˊi,$��U�N����K��B�c>]  �V��E�E#�l����_��i�&�΅�8�!06��Qt������>����M��C9-�ZY2����6]��m �*������bh����,��>'�Oz���z�$�'�"��ʣͰ�:�T�r	%8�Z���ZS�W9t}��LU�k>[s��{���|Sl?7���6�xH���cS�/���6�!����<�@����©z4.�K�����"/M�.Eᵪ����L�f�V��1����$t���rr���s���1y��'�dG�Wܿ�3�ض��b�A�jn�Y
kZ�df��p�5�6���;�fɋ�>��u�x3!��d7���)uրן�kg*�����(贵�v_�p�`�s/mg�z/�WUG�[�h4�MPh�D܀�{P�7!_��O��^�?O�W'ְD�wa��u���rvy(���y���HpbV4����ן&?G߬�a�@�&e�`�W�IG�1�u)��1��,�S
�^��`+^��%i�St�<ɸ`Pe\��|Q��7p��d hj�wi?��i��@(���y�0����g�x�5�\��V12�_�Fl,svw���D�_	�s�T�"�����7%�T�VS��v�U1�e���ϝ�Z��5+�Q�01����Z�8�H��BV�I��^��M��?�K�;��Nψ� �y���6�F����p��ʜ��-�\�
R�_��b��aퟣE��d%����q0H,~�p��K,���h�ݠ�(��A�o:N\`�8��W�Z��~����՝}�yk���(a	���@�_�7�	��g;���L՜�5es����E�6?��$S��`TwIS����GW<ϗR}ő ��L&��Y�T��4���Px}�� ��,�t�����#�o!ms``����հ�Ͳ���p�u��w�2��E��I��JL�Y��g�k����K8&����H� � ok/��,X�d���M:�(|�b׏z-�WЉ�Z;��!��T��p�DqHh���Y~c��>�r�<y��r���=�}�b?�qd�YJ�n�i�x4����U�6+T�B����_�6���/����r�#�Ut#>mWOӹg7☨6�=���"���3 ĕ����s�c�}I�N�PǞ�}��Gz�� w��1�r���H+�<�,�����kP%T|��g� ��}���bfj�{�D�$}�>�7?��=V�b:�g[�h���Y*�)@�=�exr*�څx0N�7t�j:��VH�; �│���m[�_xx��sN3b�t���$�K�Y��D���p�E[�G;zJ��@��ӌ��mZF�-�/�g�X�M��Dԯ߶���z�7?;j���N��}��as��p�^>,a8�-MX�ڲQ�,��S�:�O.U�<��p���̔\!p�C���wZg����AQ�n���Ǣ��."@��o�]�t)*�p�]ғe�.-i��?%�m����5`�!��i�F2xv{��%	��M���Aū�����3q*��e�|cl1��\��]��I�x��y�w��K��H��9�m���1�r�B��:���p!b�}-�"~b3e�����C C_
�g��/�~�i���$B�1� �M<}IsP5 � cb��7V8���׸~��g?<��^A���V�/B*��V��}�q�MyIc0À�<UD56��/-ͻF�y<��n ��HI���֙��o��z4�ᵢ�y�����)��O�p��������ǜ�����9bb�7�2���׮��!��v��J���5`�$�m��L��H��������������,Hxri�u}f1��Y����0v��z������J��9����)�%t��;�J�=w�&*�G�&���9�e���I�"�)z���y�M6�I���)�+�RI��]|QF-�rjB锗W�n�TL5_1�����9mUf`P�;=��  �D��E!�w����v����W���Cf�e"�æRV> M
���8���7 �w!���O��gFw(ߠ����5f�je �O���^�u~:ףj}����ĤR�.���4�U�s8oa�̀�zѡZ(�4�i(�_*
ܳBaAl��3�3������wP&
YV	9������M�D$0w�A5N�r}�f������zj�08QWr/D�+y�/J�����>�(	=.��puMC�d��F�=�W��v�(
�������Ks�$jj�%����bt��х�/�.Xq"��AT m�,�T6'n<|n��m��$`�S���==�ᆮJؠ݄�3ѹ��ܫ P�ֳ��BSK������<��κ{.�o�����g��O�yb;!QWt/d*T~ܽ>�8{>c���WD��h
�����&������*�����'���?pd�$�:T�\�g�YD�Z;ՕO�ȹw�k>L��&�}A9��L�	 B>:CǱ��� �
��C\�v�n��t�v5�d��OKW_x�����A5������5���YR�e�ʘ�=Y��C�|��9�d���`���Nm��Z�ݎN�H�I���C���ߋ����A�F7\/E�yB�O��p�̽e�"�٭/6	�
1{��\-�1*�w�^�ۚ���k3��]�)|U���Kڐ�G���u^�2CQar�c��?:�����X�`�՗�
������8�x�]Jl���:˜3�ޯ��]��ٽ/.�/��EWD�>O�<@Ά41��5����ݹ�-+W������.��'��>&��}V�,y�'��bDO
\L�C�D���2N�CC�� �����C%���H�X��C��7/���ߌy�ZN�͈�c3�����[����d�h��Pt��jD���>&��ϢYY]^@�}��2��"�Ί��)���O7{n�d�K�����Ј�D�B�q{A7���'�� ����s�$T�;���PR[��ş/�y�Er0�x[(MY@�"�"`��YF%6�+3L(4:*����J������o�������n���?��כk-�u�_�G�@�:r��K��F��z#A
)?,�I���&��.�t̐&U?��%��3f���1fCI��^��|���C�e2o��t8��Q�s�~���d�"NrA�8�M��䷲�T��@�ϟ�١ �M�?�H} �z �g`��)���5�H��Q�o\�o4���B ��fr}���p�޹D���@�;�:Kb5�tُ/���ۯ!؀P����G������b��.)�K�u|k�U]A�+��iv�b��h0P�L�@�|�61�'���f���R�|\h���]�BޑI�0�EԷ4�'ߞ6=��zPti|��rkF�N�����W!x��00Z�KX�x�|��N �F�#7��Bt�ܔ�<�U���U�E�_/~��mvz�Uiw����µ��XnnD�+w��f��������]]��鱬����"��j�q"����Z�hd�5��\�#�#��ƿ�q�+*��D���.>�W7��Ð�,�k�JNdu�3�S�*=���U�i��ߠ�q����2e�K����^c��f��c[�I�w��ã��њ�j5+�p�@�c��'���ȱ�hӑ	W�X�\p
:4DQQ[��F�J�A(ʴ㡫`�`�;h�f�UZ�Cg6.m�m�ͧ3>�ٱL��l����/W�;Wapi"N	�l]p<e�!�堖bwa�ݓ9'AA$`i�ﺦ���o�v�L����Aet����|��+���Ԟ�4yyEӡ�l��6�Ax�OJ,&�6�z����	26�3G�Y���NRB~�iv�z��u��}+)n�CݓaDMu�Q�~%ᢣ��D��%}���ee���&V�}�?n� �*�/�N$�T���i+�\,�J�H�.2f�XO~�L�"	^�p�J���B�L�+�����w�O/����̎R]cF�N���}�2HT���8��x�g���:}�0���"�jͿ��˶���M���%�n{]�<$B��<�KK>�f)�Y�*��]Ӹ8��L�F��|,^�'��i0Y��a����ُ
z*i��-�a-���n���6�|���fa����C@f������Z�I�#���<����ebK�+�E��ؿ ��%�4e��[~����p)c��d>�s���l�mZ@ �)K�(:1 �%�%*���M0�4:����~�;b׍G�@��Q�us%��7�ಪ��y;?�8���>žk��>K4�~,��>���Y�ε��y ����"\�A�K�Y��r簾T"�D�d�+����?)
�T�����Y5�}��MY`^D&p�UW�_%�J8�ַ6��Xھ�#"� �:1�L>�#~QRs{�h��T�wXQֵ�@���ܰ��E�<�������r��Xdۦ�/��Q�o+3푆j��7�U�ZcΕ1y�@��i5��B���h�̂c�Qr������ձHE�X?�=S��F���;n�N�@2��Y ����o�\���8�qTzeׂ���uu?e�O�F;��Pz\-l�JQ��7� �O&1n��I���/~�z�bu��玛^�	B�W�(Hрa7&Z������k��?�c����؜x��C=c����|�	�l���ˬ�kCE��3�`ڼ,��/�}��iU��p�.���-�����z
���n�^������n�.��n�����.��CBi��w�����}����9s���;s߲y��X>��ȿط��ю���s�e����\�,T��P(e�T�ރ�Ŧ6��#���1H������Ħ���e���u����	�S��Qj��*�	�7��m�Ɠ�H�ե��^u\\IBhh�$(-�Aȵ�f�Q0$0Lu�J[Gb���e�(���Y�OX(wMy���C�FQ���<\j�ޫ�
������#��g9uM�2P\�7�$���l���&8��a%Ұ9G\i!���1��4=8<M��D�sG�R.$8�t�i��?O		���{�)5�A��!i!�+|cw
W(+:d~h���'̵���X����8)�]�H,��f9C�%�c�z���CF��"V���ĊەC~�E"�Q���j�Mi�B
����ZS1j
vn����&��YHL��y�H�R�#�5�������a��8�߉���l�~�+�YT�w�?�`��;�-�[ڨ�=��[H����M��	e<p�J���I\�V�T�IN��+�G�NPʏ3�_�6��ް��&�C��4����l�;�)$�@\=z�,x70�{�d�|��즨�<lyg�D�ж�����gBi%����&4t/��-�NH��i�~?���y����.�b&��Y]T W5���B{�zGL	���`T���{����F�Wخ�9{��Ӻ���t���|���{v�e��$M�4 }d$J3v#Bxn�C�i �pG�����p)���{��3a�_���.�|]T��5
*�I�{���@��!fo��p���>���l�C�_�Ptq�P�D�Y�`�a�Du��s�����8T� ��:�	h�����\> ��/P��l�xh��s�W.L��ў�j���ޕ_m��6���+Wb=�ڰ�l_,*u3��W��C��Ζ�q�:�M��W�c��\�>�	��q��H+N��7C&
�NR�Y�������()������
ҍ�� � X)����&#^����Azr_2��_M��!_�a>ሃ��k>������Q�Im	�imD�v.��:H/�Ɠ~�m�7�Ó�$�%��Y�o���(l����p�Ψ�1m1�����n�oG��$$�aK����&�ew�o3x���ʊ��FGX�:��2�(l�j���p�1C���4�&�P+�eZ6:{�vpw8�pD�
#���P�SQJx�����G���q���͓^�3��Eo,���s�Ϩ� K�&9J�04���yJ�h-�v@���P�����TCoͨr8��%�T��c�_W�Uz`���o����O6HW�+��Н/}!��7��5h���{ 7�'E?�v�F/���K���A�ra���(a�$fx`�ġӨ�C����Of~�䄧�DG�
�R��?i����p-u���G�C�"��/6�u�X�A��\�	����  ^����-��	T�v��
_p4�<yk3a�7ü2͜��:��섕�Ge�"�l���8"w2N��|�yb��e������g���2~�6αv?k1�~<�������ƀw#6�[�E� ��F��F �Eڂ=B�@���_p��\��^�ƫ�zDǺ!�fK"�\�^��/7e�vA��WzD�,:\�����C_#jk��F#	T�QX����汃H�̉�i��2�-��n�����%��<�����O�9+a�w'�߿G�Fي�%MH�_�:��*��UT�ڄn���Ʀ�e�x�LD0�?�E�����&��5����#zf1bqf�ۥC3�-v$/۷�ùW�~wbz�^��Y�~���|#���FX����oɺ��PYH��O��6��|���6�	�DnVW��!>"^��m�9/Xg��τ&d��*��FKD��G�Y�g��#E"� ����� �#Vٓ �=�{�h �����B~��GL�1�
����*& {��@ 4��B�����:%1�`���x!�	��k�~��:���,� �M��(B�������q
0�����c���]��L�ڈ�L3! � �7��׌��ЁvY��x���7G�$��dX�@����Ƙ���]	���2�C1�\ ى��i`僀|	��(`���`,����� ��kC`?���<��_�=��8 >��?rQ �HC�9�L�_3�L4���杋�� ���@�=���SDv1v2���Ձ��F��y���|��}�O���c�ՁG�z����{>LsMD8<D7�L7(ژ�<p%�,7���p�D����fi�@֩�7��\rB�;8�J���R��U6ǇX�6M��T��&����da\�PO�#A|A�A�m�Z};�$��	���Y�;�}J�O&gI�r%���yB$۷."�X�(�c]0�(v�"�3be�1��u\����P��T��$�Y����xu���(�ڍ,sM���X�b*>O�qGv 8x[PR]��f\�`)Pg��6���el�a�򠗭��Z�(*����g{*v�ct���$y�"Ui1j����H�"���zH�'���td��oHL�#䃴9��^&@9��~쿏�NC��RG=��Y8����$�@@��m�T���%0� ���$G�^0w+aC�#$������ט`�g$�L���Ag�t۱��06��^�����֩\�0�G���R��)ZfΘC�<(��}Z20���8��i	�9�ؖY �m�����7�~Z��x��ե
s42w��B&	��J�Y8�ޙ��:��F/nǬ�2~��ᩰ5�d50�Ӥ�2���S��W�d�zش_ْW�@�����9��Yz���G�T�ғuhm�a��+�6���wB��9����20
�A�� M]����Fa�X
@�~0I�{<�۴���)��|��-X��n,���߯�0	T�4i:���)Af�{��#�LZW���;�����z�;�K�Z��y�p��R��A�1O��GK���ɹ[ۨ��%eZX.�n%+D
O<�\��F ���?�'AKIɏ]Ϟ�w	�ƢN<Uj$�����F�C���������U2e�T"���5��+Čp��y@�k\<l!�mt����_[Y�c�Ld���B��RvN����Ǒ��m{��lbIJ��&�8�\j�2���	�|��R^0��B�'�JBNG���(�.���ç_��L <� ��b�R!qh_��yD��4)!�s�(����W�G������eպ��/<\
����,.$��W���
��ݍ�rI�u���c�Tn���4�����*7�]"�W�%ͳz�������gZE��� �P�&->B%��Q����Į����9�x��=�r�:��7��M��w*	�ˑ�g5R�uEy��tk��)���%�ؾ�˘�yғX�\+��Y��? ���N0
�)f~QH���.�	bs�_��Z��2�5ս7���V��výNr�Z��h}@S���ߋNe�q�6X?NmT����m��m����ѹ��_#�v�$�U� ��~��j_��H�\0��@��"<li��ț�l�n���AZ�QRJJy$�9F��Ht,�����H���o5��kfb���2W�'x��;�1=?�0�KN��+�����c��;sXWQ	G�"��4c�����
A�,۲خ߳W�9�Uq�W;s*�XA�,v�_M��i�2�_�/�[7��v�HKKW�yy�|Kx�+Ǿdm>�k�_��z�1�D�*Ll5�>C�Q=�"�D�emP.�X��]����qǥN�<��ieE��J^ş����vn��iU��}�g|�'�ڴ��	��\��KP= ���~�Hy���1om=��$V�㝟x�t��^b�a��&(Q;3�5X��6�d_���ǣ��S������a����@��գ�n���ބ�adm�#�|��PmP�n�f��T����TXu�y�u�U����_�&ݾ~r��\Y[/�~����Uj��ū<X&|k@6���3 v�ga�[O�xz���F��3����?�2���/��u�O%W�?������0ޫ�*A�u0>�H�1ޛ�%���OnS�qMfHH�(�$�k��w2��+��7��CDȤW'5�\���ޛ����ʩUg�įo`a�F1{�r���R�
���!O2���]�v�� ;�h���꣞��ХAX����5C��q�l(��8���j��6%@� �E�US5��M�R���	�]�]0���G9q�����)�=��G��C'��N��"�[�I�A?O%֭���2Н�����糍�_YPy����v|~7�Bf����,֯_�q�|��>�Lxh��l��Pm�,��Hx'}��W\|��r�=u������:*��<5}��Z=�;O���/�:��KU��g[���7\k$�o3e��X�_�(�\MS4�q����usg��M�nGG���%x7-_�]�O�U�Zĉ���v�X�Y4��-����@�Iŧ���w��o�Ec~�'�6V�E�wE+t[�P�##qJhj��^Sm��>�i�_�e���U���J�v���F;��%�����M겧�|���3��Mh��r65���v�g��4�4���vn��kIs���'噿�t�1�=�����2�xj�ٶѲ�M}@�L�+��	6�5�-c�f.m��f{��}F���'�򢜹r����z�F�~[��������g,U6'��S�H��l��Vos����%G$�6eH|�{{ζ(9qT�H�R]�i��b��YAަ����lXϤ�2I�NѶ���QӷQ�*:���n������0F2?��>�>�!��ԿY�Q����j��3I����֑����	_��댏���5�Ŧ�ٰ��f�@��j3�|͕���rX�0�3��������Z��*o�J��i������Pi��C9j�(8z��hT4-�J'%��O�,l�;��]�`�f�()�;�f��l]��������@j5�U8�w֢���}ޡ�<~H�	�T8]]�4|�1x[�ت�fp��
����m%(͌�R�vxr����_P�!+M�5k1��s���Ό�4���EcK�Ϙ����ٸ��R��>�m���6:б$�Z�� �Rz��7�v͍��8��p�]f�}wδ,F��@��T(^}�;�/q�j�O䝮�+���`�&��D�0*m՝�E�+4f=zH�\�,1e΢qG���st~^	C1�;�q���'������e#[��ơ�w�J֩�����m�p�Y�~Z�¢��O�5*�Ҷi���b�39n��\��]2!�I"��g��q�����?Ȉ Y���&�/q[1���ϣfM7��>=%�w����]����x�5d�`�3�AtC���﫷kMM�hGɑ,z�2W�辣>��!�^��*�[���&
A2�z}[HM�]�I��������h��ao��|��՛��aC�F8�����dɈ�
u=ej]&!/��I�~j~ɬ�m,�f�B�̇�8ң��Y�6<��7/�ۭZ��v`Nc�����yQ��Q`@�ڵ~G
���e,a����O���2����D�*��4���,Xw�z#_�s���ڝ��v��;=�ӶF6��-��ua+C_�� j�'6[�z���S����~�M�'���cg�Cxwoh��P���x�&S��U�\��7��Ļ�����6{��q,%�Z)���j�C1�y��&��T��&	�M��F^�r;m%��jg�O�@��D�8^7]�~�¯�������_}f]�����)XF�p�U-V+.�d�U���6�{L�WC����8��N���w;t�v�m>��s��WV�|�>�y�m�N��Hr�1��߫9`�S���U�d#��C6d25�a���`禡Jq�[��T�f�;��]WǨi���+�a��ɡ�'YY8)c����r�R�ۉyh����=���_o3bͻ�KI�#��ݿ�g����?�Y��t.n����N���0n��[\G����UC�ۄ� ���z�".&,N�"�2&%K�ޖ���G��p\O�g��흴׾�E�@�<R�վ���Iemd[�������mY1,y&<Q�{%l|�t��V����G��F����5�l7����H�7�J�GsӶC���lDkd�q��y_@���T���?b������g1D�~��6Xq�vV5�aI΃���c�������C�d��n�n➦��n�Wn�K��;���^���ܤ�9�㜏}qK.��y������x��b��j
���J�Y	����[�ͭ�2�>�BR�)��Kҋv���B$����I�k��� %����?�qЕ���^'YӘӾ�@e�KN?�#]���ڨ��R��'����ϵL��f���J�7����ܙ�Ÿ� wL�P�7� �{��C$
yLGP��1 }��

ڈF� �/
5�Y����R�j��
���EI��;��x�'̵�xO�W_5��@�K��ymn������z&ju���-�/�Y�<|TK�3.7J���Ê�Y�$���UJ������]���ى�Q�I�+�1��o�I�p�rz�Dj�n߁�����RPk��ت'x�+�\���fo�gG������[vxʴ�O�Jc��!΃��Eu����K�ndUrR�
��Y����C�h�#����樓c��ܻ�@R��%pzn/Fܶ����=�=7��� ���!�����dU��s#�=�aA�~�הå���
��_�9'�TM��vfڲH�#���\ҶŲ��gB ������
�XP�[I>����]�E~�v����;�315)�YY�R�C���x��?���a�Μ�Z����go`��TЦ"E;c}k����p��A��5�1�Q!�Di�B�u�op�8}��=^����uO*�����{.���8��$+��{?[�]��s톇o%L�ޔW��P��"a�����)-�B���]l��V|Lq�{⟤�g��V~+>=���o6:4��t
��T(������[��R{R�8��ɻ�5OZ�8f�r��7��d�W��xb�H,4���84]��ܷ�䐃!�=;�����	^o�FL�#�5xE��x!����m������]�����IGo���s���%���n�*z�F������qo��NDG� 1BG<z�skA)N���i/%�oy����:ُf�Q�׿���2Jw��m[���J>��uD9l�F��X�ٸD���I�)j�D����C��#!�_������zؖ��HB�*Z>{��9È=��A��8/j�jc�؝���H����c��,��P���A��g��j�v��
)�l,�����+&(h~��~w�����:X\�J|�$���N�l���d*�����9iV�$q�i�⓪9)�&ڵ��9�	�ߖ+�,�4�J�4,�^��u��sf~!��o{54�ƣ�dMv>�R�$�����a�@~3�A#g�Ol-�l�~�R�Xe�3I�x���s����@�M�\8�(�:���&hH������X��<��PR*`���ӧ({ *|;S�H�H#�X�7�	_ ���mS)�-�m��āg���b�"k���g��3㧣S0�m��j8���F��~Z�h�Ż���fC��3�ë�E�$���������fo.+�'s#�ȉΥ�Ѳ#�%n9���X����2#�S�O����s=�|�j���7q&$�F��6�����w�8(�;�e���e�Z���@�r)�oo�Mrko7�g�Na����_��!�G~7��{��F(�\��or�|��z�p�Ug�T��Pdq�ט˲��e�����u~��Q��ޫ{w�G|��@w�
8L��x�����B���Ƿ�͹Zt��mu�+�_6����eĄT�4��Y(�YNpHX0�\��d��N��\��"��qk�b�n������ڈ�x����/Ls�z4"x��_�Y��D�n����aj��.����Gb��(����L�["�v��c���G��K6��!H�*FIs�������������W��Dl��1 DT�����L��z�T��=_K<,Fg�e ��
�d�td3���y���W&��|��0����o���9�YǙ�fC�ȇ��-�Û"P��NG+�O�\�u�O-@*�r�v�"�⃃;de>r�k��q�i1��jI[W���(b��xE�Zf��l�g�??;zFR��'n��pt�y�z�O��=k�AGl�U)���]'X���8Q_0}g��%����n?��:c��$Fw{X���{��یVDn���)fw�>�]��;��3��Z؝W�.��I�OɋB��M	�u��:ݖ����:.��!�MBP�]P;DI��y�ʫA؛�!I�G(*��4�ȷ�2nn6�P��P����堁Gp"&f�E� �������oE��g��9U����0�����������%� �i�ȕ� dR�p0<U�/Oi���P41�����5�7[���SL©7k؀ur��Vq��h�����e���,'C$�
�qC�?>m�T�)�`
��P���fٽMsa�Y��Fq/p��Q�չ�\P�I7�@�!�#�,�Z������|�BZ�r�M}�FΞ��{Td'��!�ԙҝk!�j3��>8Q�	Bw�nq����#��v��yjpؑq �h$]/ �L	�RЛ�M���]a�c�766��-Q��#$�]Ӳ�כ���:��O�D�*=���(lU-Z��f��P�:#����6���
����w�Y�W�f������Ê��8 ��5�ݜ[���~y�&q��  ��m�P��q�R~&��/�p ��/Z�����]�4�Q�TD. ?��~jU_ۚe�gi��ݮ�Z$j�hh`~��rkG�4d�	�)n
���-��모 �w�t�r&�gqo��<�p0d��q�S��i!��g@��	/~ՓRٺ�����f���fz��$л�m�
���|�9Aշ���OO�7�O;/&�NO'��[�c��j�����ȧJ͆�Y݌iU���:WR%^����`t?����vW���@�9{׀ϥ7����~�r؛w9L$h�C���.G�Զ��翃8�t��WT��;���ά昖�Q�a�4Й?K��lji���&�vS8`��$]�^�������/�k��}Mޯ�+�}}x`6�y��]��śY�L���
y�b�4H"=wL#yq��-�����zI�����w��)j(`^%^YM�;��k?H�#`�h^ȴ��z�Q�mL6�!�ޮ�x�6���~5���n�o�>���d-WQ��@?��[��2ş�o.��c�vB�J�k���Q����g�����3Y ��&��!���+�¦⽑1!C�2�؈ٿH!�ԄQ�Q�)���&t$�q;\�Hrl�B��\��J}X�B%2�>�H.^�������M�ڃ��Pb�2��V�ـ��fYԆ�u�]�냮C"B���N�8Q�!iTu)
r�1�Ȃ���%���`�"��V��}YP�H.�ʗ��7R?�=Φ�����^~)@���)�i��	H��moy�;aW�Ν�l@�t��`H�����5�����"2$�']JE�!�c]�.���zs,ܷ-��(X�nr��+ Y��A�M MQ0�6xYM���r�5���7�3�Pfn�=��T��y1��.�7��d�:@�{h|������8O���g#ٟ]�╡&;�x�v�-���[��)��B��gRj_ޜ�i�^!/-`	���h�вe�j��J&A���3XE��%Ƈal@��H8�6��t�YJ����Y��b�f(���,{�ό�t�)���x���:�����y-�%cz��n/2J
��2���l���4�g���$�,���a�J�G���Mޔui\f�����������?�a�����97&gi:Z=՜#��
_��]�;m��ځ�[����_�V�$.k� r?����srw8���ڲb^㊚tɋ�� ��qj�^l�yڒ���>��P:J���Yo�l�?��}1^�f�s�����;��w�� �W��*��W����ï`���m�C�����j�-_�?԰a9��@������N��i#ˁӄ�.��l[�g�^��:�n/���$έ�(hJ6n��؈��v�5a}��&"�g��9Q������)N��y#��:�y���Ȫ�����z��{����fUT���l�����:���獉x�{L�ʴ�d̔��On�c���Z7���s��N��r�	��Yǆ7�pȟP�o��-S�Y��>
���Y����& w�5�Z�~qI6|�6ے��ъR'f�1�ϊB�~R}�v!3�����N�?_o|xIm
p�0!��$���	�g�\0@S(L���1	�s�{�`B��-��^�s5��GK��f�Am���+>�?{\�d:����ل}�78�E�X<B�H�U����0yE@JJZ�٬�#�̌�M���(����P������yO��y��oK�l��2�˦5�"��b�L� ���ojh�uk߭fu�Ƣ�4������J�U�k�珙�Z��M�\Q�z-6D���za�:��W�>���N�8�_a�[�����uhE�d����m �q6-��P����'�F>1m/���?���;�b�i�fy�ۀ������^�(f�� ��{��n2������0%ox]�̙�]�ޏg��`�yv�O��~�̟k��@�|�z�.9����2���U�w버�vۚF����q������+j7+Q�-`=<�:q����7�SXpd>>�H>n�Ds�
��*�}inv=�GVB~x�I�K5L��,(e�%Ԓ`X7W�*�x���ԗ�`G^���u�J�Ro�Y�H*�.�")��k�۽Wm��Z���/�vI���-o��4���ޛ��_W2Rn�E��� ��sv�����/^E-��rȅ\��4V�s���u$�q���>~���8z�[hr2V�E�]�U��N�l��癭$��c-v�R�/���Uhl��y)bxnW�n��e.���`��L@���{'���+�T��zye���:�LT�J\��]^6�&D5��
q��?*�w�R4�WmY�o��oߟ���A� �n����M^�-���7nhw!u��
�4��7"���V{x�u�����#B����1c��G�e���+�\���!�8�.�˨�����d��֦,�j��j��>d|��1�$�T������b6����k�(u0,(�/	�MB��N����T3���h�u�CB�g�˞9�B�'K��l9N�$�M����b������Z�ga���*��b�HH��4��@gͧ�ݏ��n^Ϋ$�%~��U�Ȁ�����X�4�i6?B(��Zu�8��Rw��'#��߆�L��Y�i�閍;QR�6s|�)́9$� ��B��q<_��#��|a\�#����Q	\$N��=j^����H��z�Mrˀ�y�Z�V�C��QeU�2�Sz���#"���s��i�2;�e�w��e�^��">�8h�62�̅�%X�?޼�V��Q�=]i��]o�=�S�gI�/c�oX�q"Ǻ�mr.�/�rq���>�s�ػ[9�_���)[m�rg^bURiE�Km)r�S�Jn�9f:*!2HÆyf�N�S8�X;��j�)]e�S��Hz���g�[^t�#X�tq�9�Y�q�p�s�����U��y��J2�n`j����c5e"�"�n`����>�R�����\��tg-&QՋ�6��V|����������t�b4Z�f���$�����"<8���8E�$���0�l�mڧ�#|b�*>qV/�����f����J�u���.�����D�<�7$�D��<��t6�+���T�9�8�6�'�������"�f�ń|ؿ�,ȷz'�Ũ��3#�����k"��b�%���xN����n��-�lL��&�[fg)Q��K�4tBc�ִ���{B,��5O���͟��X�6��U�-�����<������ރ,m��I4(�GX����󡤊d�-t�8&
W�o�M�y΂B_Ү��.dYZSd���d�׵����rF(3o7�����WS��x���O/˚X��ұ3�����TA��B�u�?��>�]��(0$�y:l>�	*(���v�a�t$�v}B� ��x�!�v�΀��Nm�w�7�={�}���v�n�m�	�#r#�y��`P���}&���Ԭ/����u!,HRlX?�y�h|��\�h�1�w�֍!EAN"uv���]��C�y��$r�~0z:G���<nD���|n$�CՋ�&�r�Nԝ���8��yP4��<A�❎_W苾��7��Ⱦ�����?c���gz|j���ɲ����!D�d-���.�hF��x7�󡯹GJ84uF�ɥM)Lbj�-!�B�ǈ��8V�ܿ��%3���=6�O��x3�⵿D��ў/�1�Agd�EDm�8�f�/�޾����OE5��o�}�adv�ԗ�斾��'�D�v�VɴH�"��"-��s�kܘ~x����X�#�"}d.Y�;Dx󼤕m�-�_�n�GK��x��������߶��&H�{{�4�k�j4�pr�Է�-A��>����{������oÜ���x�G��2c1����p��4�]Ь����`��]T���z��~�fQg�(e�x6�M��I�=hgH(�]�'�?f���=.�[�H�g��/�h�)�,�|1I�6�d	L��!�zt�������@��Mh��ʟc��ҵ�m[�s�SH����|��f� q�d�pU�~�w�r����w3�e��YI��R�r�=ٱDH���kC��Fl��y�w���3]���B`M�����h���#�E��H������n8��`퐲
�K�n�EU��5ii\0�$��%�Md��Ekl���!<�E��1��[޻�iB�)�e�t�}�������{S�@��0��0�d�yQj�S���䟃01��m�K��U)\sB��ŦMxBG0�1
H���&J	>�q�f[P�f1���@1QrX��2����գ��Q��O�D���s\���L!j5'�Y�D`����g� �0�8l;��
"��96�)�A�x2d:)Da��R�,c�{Q���JJJ�@�',E�$��̚$P�c��t�^��T�2�%%���c �B�sCxE7�?1������YD#PL���|���>���͠% ��'�GH!z$A��_�L \F��@q	�Å��B��,���i$�OC�� ��A l��DY��� ��1dL=v�)UȘ�a�7�Gm�cF�멂B�2&��y���<d��;��� hMA�cԐ��@O~@$���(�_ � # �2?��	� \ ��Lq�z�\l���	��-�ƀ���`˷@hH���ɮ�TK A����_�V����d���qBHH�����^�
Ї�	�U�7��� �4B�O|e���} nVA�G]".7B�&� n8E�`��-NY��9�"ȍR�jV�Y�X04�/
w�B0��C���� W��}k}���G.LKu������J��ݚJZ����\�Aue�\D;j���ҍ�n,}�He��
�su]P�����R�֒�y�z����K4D; f�hp2f�U���n�J(��t���!�ȡ�ЬGXE���a<��|>kŏW���%�Wt 8Z�� =J"�%�ݖe
�֢ʐ������@�]��z�p�}�9W�<�II{���eL�:p�)�Yc�z�)o8�PL+顇���>�ô���j���������3<�0�1X�#=��q� <���ML+�����a����ĢD�oH��F���u=���@�A���ւ�B%����p��С�N_��Q��ç~���MAe)z\H�T�Ѫ�|W��LA�2h�ܲAl0���;1�nO��%������z�0����RZ���C�d�Jf�O�[5�����.y� 0�̓������. u�OH���ej����#��J�<w��&%>X"њ�{��f�.�%A��H�׃5&$�2M�K���	M�
�#��Ats�Ε������=Е:�+�E�"D@�����YDm�����u�"}�~nyv�VZ1� �$�VLF&�2�R�6</�Ĺ��?�CaN'��}G�̈́����CH+�m�+�X�9����`��\I-���n�C?���B��p��s��Fɰ��'��������ԗ{��=��j�Ik��%3J�mw�]I�bO6���C�V��&B�� Z0��6{���|c$�4%l���=#�2	�9�F@]#,KQ4a��A�[�����x�;��Sk���䖂�Z�T5�u����[)"��2v��wA����[����?P`3J(㨈H%99Bz_��\����b�,�v"L?��D(L]$T��^H��0�a(�55�0����J�JN�8Jəz�!���Mͺ�Q�!۫u�4?�k�� F�%,���,	���/8})N�o2Wc�eպ��̷o�۪)�NK�wte������d����3��R@�i�:ޝ���z�TdrX��Z(�Bd��g��	���P޸=�:`�Y_0�!BOa��X��Hsr�z�)�u
,��(0/-)�v�z|�v��]d1�ߥg�i������ć�דɝ�
tb뜾�%�v���<����zT���PW}	�3�,�{hx/�=��$D�׼�<�z$"�Ӫ��.��`.����2�&���K���C���Nw�2�m�J+_n�%
dͽ��J�φ�)y1g�������:�m"�b'�L�pU҄���@���7��w8�� �0`P��(�����m,����>sl��;�ii�Hʭk�FKNr80ڜ3`�;{�E��s���i9��~^آ�GC9p�?�r7���#�
���I��K�i~[��4,�����0��`9}`���c���eE?�a9O#W�Y� =�f��с�-U������M��@��z�G������8���.F�?$ӿs�C�/��ԉ�6�j@�V[;�����	�A/(�O)/�B޻��+0'��u%8lG�`70vk}G
͂gi�%=��B^q<Yn�����'\Ee���םߴ�:�ۜ ������.C�^ڣ��k�tf�B���<s�n�W������ܻ[��n�͏c(�\푩{��]��zm�ٷ�6W��w{�y:���УPJJ. �����RV�g���У����̛�O�]CԳ"�vO��?���`�� �3=%I����@ޭ�D�uE&�����o\?W��=�ʳ���My�z��3����4K���g_ֿ=t��i��7��j��
v���������w��0����F�Ni9V�N�ibF7	��h�=[��~��M��z�tzZwv�����Q���dK�z(�l"`<p3�+�y2��_Z�����e�&j� �"�t�9W�\c�c���"��-�Xi�F��Vp_ֳ�\��rdL�r����;.��7�0S'�DO��E.
���EW���zsa\�����OnE��J�*#
�*8���B���DU�Ye�[Rum�FS�v;�Ы��
s۽�|�^��/�YIH+1]���5���Un'�+_/��U�	������|�K��rr��Vh1��VQ�f�D�Ƶo�6�x[︓�x��#"��5o����ѓ4��I�(�	lc�|&�����x���m�׹���c���S��8ΟK���{C�^iԹ��\a�����WN`��<|���&}��ix��(_}��*%}w�\ܳ��'X�J�h��R^�:�k�뼞�E����wk�ظU���x7��sy#�	]4.�V��t�G&�?0���㥿�7�;�8��R}<�(�&��;BMh(��A�K\Ҍ�x��B�:�5����d3Ld��U����w	^��H���>^v�v'i�}q"�sSl���Q�����t戻`��
+�����㺂��j��Dna�ͪ��D$Y�l�E�o(\&���a�\�?CJ���	+*��頱7�"~<|��:���o�'x�ƭ��ة���>?P�i�V��9��uP��ww5l ���6��"��1�r���Ź�����3�R��V��u}
��<&²(\@K�_L�>��2�I\wҶj�Ĺ�J
��#탡gSBjF�ƒ��
k���#���7�x�����FOQ���g
�?���:ck4��������Fz��o)�1;-;���*�[��?5 ���Mit\d���Ģ⇗�д��_<��+Q�ZQ64��Mւ��e�R��W�*���?^�^��DP�E",�̭.��u;���R�U��
?F�AVn4u?f�����^������>�P�_F���/��q�d�m�4�,��h��{qy�˾y�h�IP�?m~J|"y;p��$�R���F2�h���%��ػ�}����-EG� �E?��l�	���M�C��΄,yL��4�g���}��5�8�?C��.��p��٫4�mQW��,��
=	�һ6�e��H���x,g�:���.fs��@J�(���8\ǷĆT`h��n����t�w��f]��6��@�������$��,����}I,����j���66�P���k]{i�y�oI\��*&��Hd�O�Q�:&�D������7���YC(R���
Fwy���1=v4V�|˪����������i֋�Cpw'wנ	��N� ��[p]48�eC�8���w�9��StwuM�SO�T�HHĊ�IdE@H�Y,��[\�� ��o1�x�U�AxÜ$��i�݂V�%��SC�	"`t��e���9�D�x����!��F�d�������8smK�XWE����5Ua��i��Q��K�4���x��qS�Y�q󩡀�XP��Z�V>`]@}��Dx��D��v� ��l4P(po�o� �x�6ɁE�����{y�<jZ����mxR�-n����������*�rg��(��V�y^(<q���J��h��u[�,��V��ŗ_(=�hv�d���r����7�%0rW\�~��72jʱX�f� ����].*�m�2Э߉���s����:�����3��<W�#dsDX��⌬(Y}�[�6,xb�NM�%�̻첎���jyJ�]�2�iw��|l�hx�\�s�ò��b��45��9�*�p7ћ�yR��U衭��C��<&5_��)�	��x���rb���{s^�u��Y�ga�F�u[*Cr!�r��� h'tK��R*H��go�t��V�E�z�ѓF��=�7�w�R���o�UٌzL^�?��K��(n���;:�\i�4"t-�4x5֑_|��MX<�׿`Մ�}�G{"�r˶��������z��2q�^���?��f���|��G���Sr�s��&_����d�Z��2�_��]� &��w*Z�r%[s���a��(}�Z��gVF˦I��ܲ:���#�Z'>����dv�w�)��]��	�)tb�<+Րe�=�vվI���妎b���H�<v�7����/�z<:Q�?�q��M:]����u���ʴ�T��΅MR �<2v�/�J�@8��]D:�Q��%2gh�:}�,�i��9���o�/!�dwYV���^q�
�Ԋ-�m�&dl��r����뉤�*�U��6�b�M��]�y�1=�$�b����t�w��I��c�ȤR�C_�`_�ٖ�O�=yqa?޵��)�q��9����6X�|,ϸ�'0X2ϴ��H��2{�V���(��3$��s�*��/�q��#U?��@�ɋՃs�'C��/}�6���{��F�G�ۏ�\���i֡�Xb��{H����|���k%}�֝,7��`��-dI�-z'�8�:am���zE�Ǥ1�hڹ4'\7���+U^}�j�r��@*$����n$P�N�-�!p�ϩ®��l����r�Ѡ��r���@?�C�x�C{��v��K"��^G��N�WN݀�������51H�K��K�����e\i�NǺC o;�/�d�u����%/������(�r;��`���//���c�A1J��/n��P#."��h��~�H��"N4\veÆZl̘���!�� m�4,��K�j�G�iR!����۫=�'u�`'��&kt])mM�Fz��9��'W:�OB5?�����ƿ���ǘ��3.����������n*q|ij�fp�w#��*NC$�v��g�>�i�����_��<xT�t ��<K%�6��&�ƥ>FW�9 ѢЋ"�f�|Vwx�ơa�h��j����l`����[u5�<�R{3�-+������!�����)J/}���02.� �4���m��h��ލ���J�|Q�aw3�u�K���ɠ��\��կ� ّxPIG�PF�U�jd�,��rļ|��C?��í�צ�i��H����+p�џ̂�����#+T�
��N�z_���U/���#,��dQ��@��Kd��Ih��8�	��
��#w���2���H���x􍖟u�9BPCC4u����ۡ���B����1����n�{�Ȋ} �J ��L��eE�'RȖh"�/˙@owp�=��[��c]V����휾�V�R*���~��Y��S�]v��k;���e��*z��h�̞7�!&���X�Y^�	u��KP_�Y��0P�7@z��$�oC8���ғz&7RW=� �F|ƾ@�\>zq7q�J�b�dtՌ��](K�m/�����G!Z��U|�.�>��(}��~����
�)wp3H�2l��F����x>T�����5�<DJliYm�So�̭H�" ۦ:�j��t$�a���$V�Q'������|8���5���$����g����m���W3�XBlы;���O�庋�(C��H ���"�;�8������{ON�Y{��v�{�ͨ�
��P9)a �B"aO;%6ؾF�I���ʷ,�.s[��ǚBb2Q_�J �����[&���-�?=JP�/Z����o4��~_�(/����;b�L�U����I�ʝ"R�{"��d� �'ר��� �V���[e*W|P�eQ�ѩDve ��>=�!���m1��bd%R���a�����(�_ZI���?qб1E�d�.���Q��Z캨o�`NQ�NX���)A�l�w"H�Z���b��A�[��k���n�Z-��|4��
���,h��h3���&�j��|�������o��@Y�RqH�2葺�����}��`�c��-տ�Ge�n:�H����e��"�V�%J:J��B�=��i6�*"�7B�ą������6bg�6D��.��*rn��!��Х;bI!Գ�����B�X��jK3ʊ@���O,�)��/}(�7

��,�6�Za��Ҷ��7�E٭����k��Gm@\tZT�_���%F���┯��^%w�'��B���2�g�!�3���[Y5���a(1`��Ƕ��~`�uG�@���Q7!Ͻ���g"+z������F����I�?����T�P^B�G�A�W�����9����~��DcΩqB�O��z�w&:ss�d� ®z�t��3����Rm�ҽ��w�����nr��hy�"2B��Ӷ���ِtRR�mv�+�tY'�_=7L;�	vh��N��!��+�:X��'A���;���..�W(�j�5�Z1c��t��v�%�p�Ә�M��#��\@�|���/rW'��f�F,�[{�Ȳ�~���r����6Q�x윗�(�KPV�;TbJ�<$��jW�]X ֈ7�X��������,�R?N%C����E�`R
�܌���ju��	� �i�;Mo
V[�j�C��DS�@�+D �9�꿛�eN��n���q��_sI1�4+8����\��t
�x~��hyd���3�L�wE�l� S�1#q��"��������P�bd=���Q��;N1(�-�2_����b:
47��v[�;\��b�^��&�*;6]��{k^z�qл���]������{P��ǥ4)J�w܇�TS8&�ʴ����e*_O����4�N���΀%+�7z�)J��Y�ĨP �Q�X�����Y�7�c�\5d/�&9z_��b���	�of��p�O���O�9)�Id���1����(��{�ח#E��Of)F_.?���t�҅�c�"�t��{B�H�q�[�4+"#E��;���h�l-Ռ뚮��o�sM%ay�Q	�O_�~�oƄZ�
]!����!��[��z�*o�m�z����0��hL��V���_�yU9 D���ߧ�_�Ї׍���ޜL��Gα�[�>�˲o��HyC}�k}5��zuB!����rQ_�AR�wOY�26}�;�B�c)��������K,��0�3�̇���>�=��h��t�s�A����,	�u�<e"�l8��*����rP@�ظL*�y�X�,P}��mCF��^R�Y���x�j]��x>ˇ��wn%��l�ޛ�bq�4�[�����Z����~~*ri����{�7|�!�~�)�m~(���6��]�eHS�S� 4�-6�����V�E����.����5�+r��R~���1�9��lF�(Q�1��?��J� �IF�tJ�O�Jz�oO�ǡ�c7���r��P��B*��60�v��86��*`�J(�����T��y�S��@��y�m%As�i#��>��\�84z���:��ڷ̯�[����R����U�Uk+���ͫ��,`�g�"!/rF��.�u#���DYY^�?��ӱ�K�?k�� 4�D�=J�_���+�|Cy��{D9D�?��-���tQΗ���É�1������LQ�%z�K���OTWW_��tM�8�"��T��^{ۘ���ϥ�p�j���[D��y��@�_!HD=�B�ᯁ�)t��_C�V<��V{��dr�H�q���vλ<	~����epK�t0��INN/�Ȓ�{�7{d(b�}�]e��;��(�33��j�(�~2�����V�f�+rk�ާ7�'+2�����b�Ic��R..G��y�ngG"XKR75�p�ku�����&(��qSJW����ɚ�1M���Z�	���'X����{o��ߔm2�$��B��F������o_�A����x/���˟3�䥧Ӊ�>��r���@gBkΐ&���,�d~,&+xP<�5�ʹx�n������p�i܀�X�n���Yz�K')�(U0�����\�J����_�J=�Ʉ,їǕ�#�J"�N]j���L�����|����?Zdu�H*�U��{[8y`V�~
����a�y�Ƕ��(H;9�7�堣����YH�� .� ������S����ղi�W|O�8F���_l!���U�L ���b��i���b[_���Ͷtʻ�R������B%(�mn��I����c��ؚ�[,EZ����cf�>��SRRr�U�.�3q�'E>ί��=���U0��J}"��x�U\�?T�A�M��j׌����o7ye��q|�n�ئR�6��[[�|k�>���}��_�5�K�N�u�v���\V�'W)��5�x+�����^�L����:v~~�$�c�+����B�]�l�mN��}+u�wm"�n��b���qy�Gy!��o���Џ���Շ3p��8�@ɯ*P��q�@2,����f�-�݌u�� ���O���X�`]V��n��O�\��A��c�ҴV�1p��_�/G������xq��`҉��"'1J��r�~��D��C����B���)Uq!�


��?�X2����$z���^�o��"@���Z�/�>lhH"�Y��Y���x6"�y����v�W������'fi���g��m�<��S�8��7�̕�dv;/��c�����}�E6�'�@)�Uw=�;c�*�&��2����� 
��A;�nLʆ��`
�ϛh�������$TT�g�+'�*7�P�H�3����E�<0�#�'B"����=��sN4��fah�Og� ��/����c����:�;��綵�m(��梸wz����Mπ�Q��������������+rr"@��5����ɏ�b���e>����Nc����!	g�2m�:������"�J?�g�%�`�x!�A�÷821s-W��y���>Ƴ'��&�=]�:��f������'hb�l2x�FSs~x��$��V����&W:�֙$��~�E����#q��bv����x����Q>c��m69k�;?z�ld��,ž{~�L���C��)J/�v��a9]�Y��§*m�!u�z0TI$/����!����廁���"8�ը���;�$r�/�!�L��i�8҄�v�Z�!�XKk	�(���"y
l�4�����t��)J����X��P�"xo�iD��͸���h����djf����C9�.����3�}��c��j67�OJ �Z9�!	�H��,X��R������]0A�͙sjt}
K�b���L::\I�4$�*�ڒrwԛA�X�OX��z��Uâ���L9��Li^��Gg	��f�M������XŹ����CJ��ě	6Ĵ�	|:��;���� �c�oht1r����Gw�;��z�+�\�l��H$ܦ�ʬ$H6����<��Y�F�i�+{x������q�5��-�:��>M�J��	�'���Qw�"d�J_��&�����p*�6����u����W�{���)ծ�x9�-Q��U��m��o�k��#�\7]J2��hD�eD�����?��ֽ���C��X�������.���:�;l��}�dU2Ǉ[��oRA��;����\")��`��%4�B�;-�mΙw+Y��B��ze��\�p������H�c+�M���l�u"��Ȼ����w-���N�K��d�_�}k�Ά,!c��`�Q�V�KM�	g�]�.���~�^h��7V����n��z�馁f:�8���v���Z�Owr��{d{�J����Mƕ�G5�����6�s#�U����D�������8�k��8&�p�KWzcޔ�f/��\*[*.ʺԅF6U���ɛ�]�7���u�VD4
O��3���0v�]dh�g�|B׍D�c&�pv�M��đ�u��8@\A��Mb��S$Q��th��AJk���b�E�{�5�2�]����0DZ7�|������z���ߏ(�¶r�D�7��!0���F.���bs�8A��#ѯ��_��
�x��p&V��0�ND"QD���N#�ۏZ"�ʋL(ڷՏ9!V������$�@�q�<bһ�.�_�;R�l�$n���Է��qbuqq�`|z>��a/"��$�p{��#�1H���?��mp}��������v84 ��u5˚�OSiG]����_��eR��;��Y�X0oM��*�6>�U;�뷁��e��b��J���-�k�Zڶ Y,^y���ɫ�A��yL� ���_�߮��vbu;t��,�ݬN}Y������K���ak]�F����fj�A��Q��Nv?�ޓ���_(캗_��+��dmt��b����)>�~�$.r輫*��z]݉������)aˉ�X�)Z�ɣ�s�dc��E��5è�\��?QVģ<��-%�RsM��*^ybȸ9e��U�ü6W�c�D�w������<c���ڄ�$T��������s��C��!�� O�7�y�(m������ZX9k�>���v~�P<:�Vz�B��Z6�r�ȍ��~1". U�M�d19�l���\l7�KRn;�:�f����O'��9%:�&=�;[Y��vd��{n��~$®���x;	s���7q`��؉V��0Q�m�gu�^���?1�5h�ʢa�_��։�Ly�9;ǰ���!����i���^}h�pq2,m"�ɮ7���+������Epں�e�"܀��j{�PC���J>�oz�0X��]8������R�|J��n+r4��F��b>�qgk���k����Ã���@�|�Lx�PB
�wv�iQ�F&D�!p����L��t��U��i�U~h,'@���4��)�x�A�G��E������UV�{9җ��H�~����u�$@ko14�!jY_a�p��ZI*l!־�D��ؠ/f��� �Wg�V"���`�/��j�kz��`�a���
�G�s0p���'â�řR��o"�{��I��)�؇ u�_�Vt=c���?��2߂1��F�D�;&$C���䴻B���(�9�n&)�xs�#9�����?{Oh="_`9f��{"�=E򕇝)g	&������q�|[���{B�wo�/��2�Tžz���< �VF�$�5�.��a|�%e�q�,��Б�i�iB��Z6���5(YKV�����U�׹(À��,�xP+���Z	�q��g���d���T��T2��� �P��X�Tl�Qh�S��%l#�vZ
�u��h*�Jb��X��i~�T��)��G�����{��ϗ�Ϻ#�3�y��*V�ޮo>��T?�p�;��B�q�U�)Y*����9A�����	Ů(dL|��Sr�[���A�G�⛀��&�/���7:��	�*�34��G��*��L�d2���dɘ��p|���ld����Z��{��i�e,���C�2��@<"2T���/XA-_IB"]��k:	��,��)L�&��
�`�$FF2r60\ƄΓ��Kg�O"c_5D�� T��,�ʩu��*Б���E���h,蚜��yp�Xa
1�І�(^:l�f�J�0�L� b��"0�%L9o9 ]1��	��}�9���
tM]蚭�yBp�Ԡ���������[�	���*�Ua�:ѯ���F��D���7�-t�tm��C}`Cx�5�`��-j�E%��HǀjD�Hf�\آY�2��U�#��g�NK�CǦ�G��( f"Oؚ��#qÄv0!t���1��U
�֚*4D��/�*ĀY^U��Y�(��ǍT��b�B k5.\�'845��kvLv��W>����}���Մ�°Vl\NN���x�̆�!Z{�86�Pl,)�e9><��"�"h���p��#D�>��/���uR���Lv��?�Ċm�ɚ�,��JDφ�;���~+��=:>��_���N�*���?T*Ygr}?i��{�E��vme�:T�L��Ǝ/��a��U	��?������P��k��h�P�8T����Ăr>��b��p�T4N�"Ƥ�q~��7Xj%��Hx��%�퐙@�՚k������'vBK�R��6{\��I��q�H�lh�=xı��E4M�+䉛4�,yÝ�
n�#{��"�1��ό�9R)�\��X �j>��i�F0.��9�$J�S:�m��.��n�)�@�}�N�\�ԗV��J1��	)�N ����:K ���s�	]~��/�Jk7�t*�<�
!RBQܲ ��uvb �����;����OLF")�S�M��$��U�,=(�i�_�`�%W�+� �سy���Xٚ~{~�,�vI�<�=@�.⊆	��)���ЯLC�~qi��ǡ�C ����p�K��i���W�)��;���<��8['����C��%t��N-��zMm#��϶Q��MH��2��T<�α�И��Hs�}�	;8q9w�~����ާ<v�����QW�@(�N�w�<M�	Z@����!��l�_�@ri2x(��H�L��ڨ�$$[/��cg��	=��'| �͗����]���8�}�d���y���&>�!F�)�NN'Ԟ ��î��G�R�~�z֘"N:6���6>X�����v�:}
K��������*�D��Bʙƞ�^_��Cz�>�q~���䙄�^��>�ʵ�_Ez� ���z� �P?,2�{O�_혭������70���	7���ށͲ	ox(��;~�� �ꨥ�FQ$Ik��9�~�Җ����% ���;(�a=�Ҽ��0�ɍ�M�����u�[x��<f��])(~�rM*Ǹ�W�2M@��S�G���}P�L�o�+,w%�mu�^
�:c�4��ဏ�?tx�P�J0�v�_v�GD��;���7�x̎]�=�=�>H���[ͺJ�m��
Q��e`!�|�쌍W��H���F��B8�n�Ф�74+m�Y,�'}Z�70
$�6��O�C[�ͤ��r<���A����]�o�9��m��՘'����4�5$j�<�JE��c[J5�M9�oId~b Q���QE�֜]̈́�~-��o��\T]�6�1͕Z[q�b�$�"�=�rw�%"o��P�d]=�עr�~jv]7�i��3Ncr�ӡ&`?2��;�d����h��*W M��a�,Ǩ��om-� �m]��N�!� ;��=��£ܮP�h���� x�p��b�߁��j+��C��+�	�{nP�}(?�Wc��(�e�ɈEL��~��C����1����v��Sf��;u,x��Q?�/�]Q��r�GFPEQ��4R�	5"��	��-�?5TlP������#�G`A�|� 1��P?�w��&o�����@��4�&�5��w����d���K���7�]r��C��?n��w@y=mN'�`o�F��I2ॺv��d�ȁ�O-��\�!,`�GΆ
��v2�㈡�@KE��F���J(B[�\>cTi�R7PR�M��b�U1��bj
]..+�o���Ϸe�W�����z�?YA�Q��i۱��E.�\���1�����G5�+��f$��p�������m�b�����:'���~%%0�Gc��m'|���?W�BL��ʥ����9�v��;�l]���q޷������~�ތ?NO���V�Cى�|�{Z#�e�*{!g&`-u��SI�}M�[�����p	(��d:�wVds�C��%�s��QT;�>H�o������ �^�A���&%��{u5:�LD�)W��Q�K��i�1;���yV-w��&����|�j��J�%��fcM�A(�W/��A&!74��L���޿J�m��^�2�ͳhǢ�O~���{[�(��f�0�.k���ez������e�+�Q��
���Ϫ8���+Ø�G�MNn�Cdyo "�-o�b�ܰuI���u��"L	>s�pI��R6�6��!T-�r'��G�(��ZQ�%3	�vi�li�~|���/v����~I.�*<�r6X�+�s���,Y�v�cȘj%�7g�*"��CG�#��(����@����-�jq�X�ޛң���-���ȷ�.%6���n'P����я~�$�,yM�}�X@� z�s��k?�-C&{ �^QÚb����`wn�|�QN��o߉�u�$�T5�IY"�Q���Mc�}o�W[�`�?��ސm%����h�-�]��hdEt��~K�$��vx��+֎�w+�ް��4��tJ�+��Str���t�F�y�q���C#6rT�@�J�ş$��mΣ�6��>�L�S�D��Q@��9�U�$@�-�v�cJC,*u���fۧg3
�(��;�.Ń>��z���$�x�gW���[9Ky��1f��o�{���b~����;��%	��X=���Ka<N��D�.h��#���y�ļ����^�I���g�ׅ��*�@�_äg�I��`D��k'OZT	�@�t�rSaSX�;ė�<@���$g�"����C?~�5&��ڣ��V<%��e+��̳.��P#xY��F��(�_�˰�uBFi��j6B�?�6��'�?@
�����91���Q?(_��x^�S�I��:��b%_����;�6Xٲ_I�z�֢���~�w7�����r���~��5�K����}$*$��>�D�ǽ6z&7� ݙ���(e�~�b�M�)�����?��Xi��-��R����	�ݱ�5K5��*=�~��DdCV����1�9�a�f_�[
���4醗}΋d������h��,�Ơ5�"鍻'��X��������.�DG'R["�aҰ]���P�JF�^�Z�׆�З6��5�jrW`%�#h͒m2w6;��+0��<�	Ѵ�k��|�<9>��H#�hi�ٻ�@�{9e#���z��%T�����4K"��hn6���#���t�� ���ӓz!qPNy>z�'Ⴤ�VR�}6�!s����j,;�Xa�wZ2"eqH�R�SJ���Go�	}͉n�������))h{����k2���Ȱ��.{�'�峨��j����C�ى�r�o.G\��I�8��,�^���	I�o�?>e��ڹ_g�}3�ew�����p}=��i�w=�XJA}�iK���=!]�
��6TO����e��e���p_�yz��?���p��� l�m��N��|ο%���3��U�����Z�n3F/�Qy٫�.a��Uki=�+Ccp����	�*D���	T���R����	�I�F>[��OF�����:S� �#	IRj~��f�Hn���UAm�G�r֜�clT��Ɣ���7U$�sא�l���ܾ�r�Sk�$���� ���M;`�N����J���%�w!H��'}��(-��L �f�yG���}UTR��Y��r�h�������C]��V��)bA��
Ηy��Do��(�a5:�_牤Ə�|����L{�c�z���h B��Jv`�E��Õwv�(O8!��6��S�>���0�F��T�P%�w����>�TH���.��*_�����}�����fZ��Y몬۴i=��y�$�-����� e%%W�{/��Mw�N�������������$����6��K��"��%�U�TD[�M�~_�QIΫ�(,��m�冱����T*���ŵBq�A+�%ǑZ�g�sF�v��"������h�_�X@(���[�vj�|y���uH'}��E��{-�zv��]�q� �������_ח�4گ,�1�����@�{v��K���D ���/�Y����A������x�l�oF�����3lE1G"�t��C���%�/�k�Õ] Xכ�'p��?�忤����/|�yڃ.�8�lĨ6��).�#!�p)&-�`<�cS�&h��r�*�3m�ʵ������D��WD�1:��`����[[�̟=��-��Q�)�p�����Kbrq�!F��>�m��(>|?!%'��B��(��b����>7v$�B�3Yu�����Ž�ǘ��F�n�U�Q:Z�{��fM���6���W�y�0���u���{���ұ#�������{��w��B�Irj���Ht�Q,]�x��AE��9����?d̈́�h��s�@S$\i���P����C�g�Y���K��~�=;-y��u1��^�~{
�2D@���4{\�|��x��Nl���3�u�:Z������"M�h������̷Qև8V���C�ҥ�3�����N8�{�L��2�G���*p}#��S��|cmٕ�oS`O�1��Q��l�6�R��A,-�
�:��{����+'�!��~�3�4�W��/bf�*( ��Ջ���$��V��[O�i��Z<b�*B���r��6�᥆�+��7Û,I�cbb�oI��߈l� ����g��m'^FO���oty����ˍ5i�s��$7�3��JFX�l!�쪹&�A-��-�p_��:�y�d��hE/�V�f��VCx�����2����4	ȫKƸ�9aUD�U�mRi;|��Iji��}���o�XaoINq����'t�*�	!��I���	2��Y(��U�w�3^��=n��y���;�X�GW��i�?��֦�B��z�J�>��9@z�~�y�����׿���s��N%8TZpLhrS�n�7ם~��7w^�Jbnf+��f��f��˥5���"�qk���"md�(�VKeнф5/ԗ:?���G��M H�\׷�O{�B��o'6v�ǢCVZō1�#�.�O<l�8�9������
�'���wD�O�T����m�G������#�XD��m/���垆�Ӎ�����Ƞ�~d�	!�^��}>D��K����m�Qq�1�Į��K�6���AD�Y��}��'v�m�'˝�/SE��M�Hi��S���!���{'{�L��7��r/����r��7���׫����#�	��0s%jD�O'��1\)�Vfj��&��9� ?�o�/�wS�c����g&B_����&�;J�^������|
���G����ή�>XS����g.��2���|�GJH/�e��CJY#ğ3&y���Y�IzR�������1�ػ#���E-���a6#�,�拾�0zU�0�� 3���X~��s��O�2�I�� �!�O�|n@̢�����Ɂ��?�=�����r�p���+��H�U؂�-&��!l�.�j	�o��H��~cƟ1�'�i2�-T&d4�4ӷ�Ѥ�R���ƭ=��������]��E@X��2Fn�V���VІ������i�Vv\�x)n�ζ���g}`���p��{�bחʶ������HA�35~�E���dD�]��R�#� .��aa&���Ɠ$��!�c�h]*"��EJ�[Z���ׄ�lK�57�݊3�Ņ_�hDXPII���{U7>=�ou��/�+�LLVjӉhԬE>�����R��x��\>,Ҭݨ���A7�����E����8̛�Re��1��\~�W�U�\�a�
��^o�ri(p�_ř(jݜ��/~]4>��;�BS�z���(�I���W��S=Z'�r�kQd�uhE�l�M��j��>�Q�&|�_����l��,�s����"��v/8�no��I�E�W[�]�Mq�˄*0���v��v���eһ�}K!�we��Q�I3�E�1�W��%D���/5S<���k�o�H��#zi�(�Jʎ.��u�'�W�/@�6�jq!-93����������G��Gn��D̘�6rE*Wtj#5�`d�OE���P�/�� �����	U(��BRv���Ф<�+�e$	w}϶�IUGHSO�K �ʐo &�Fal�0��{��d1n���/}����C�#3j�3B�q�Y�"�YhP���4p��ګ5���D�c`�훏T��eچ&k�]礜��wa!���^���4�+E]kj_�M�.$�8�☊j��ybm��4e�e��o�����c_v/|5�)��M5����~�]A�����M��r���}�M�ܹ�eA�>���Y�MB�{��!�8����sh�˕u��2�<I�/%W��P�^�:d�#� s�H�,8����)@��g���r�q����c��
-�A8?�#��5(�O�U~4B��p�i/�-�C��焤;�5o7Y(.��eXc�1vޟ��x��Pa��'��4��%�y�0��Q�����bFkS{����i�2Ϫ+˦��Ĩp�g ��])�t[���!������H�)��� Ԁ�yI��N���ǒ�Ui���u8R�X�����n}���S�DŤ�L3�f5��wX8��_{~�G'�0�s)��|�% b(PoJW1Fj�_8��=�d���0�Iu���ݚ�H��)��Ϝ��wP,76�]�?n��N^,<"#Q�7�4����+�岅J,j��nl����U&����$�=a��\%%)>�'�d�KG�{S��$���ʌ*�$[M_W��[0f�T��WC�P'�!]g��mi"����[H�~7b�0�����5q���}C�7s=�Ֆ�ڟy�Dն��]#�"3�""��p�7��b%
G�l���RM�6���{���Y�O�=>��u�9�+�1�����aAQfJ��aJ�����_ ZEF�ד��.!��K���/��r��O����U.�NqI��6�;�t;�땻��%c�0��>̝�2�2<Cݨ�G1���јS��C�<5�E�(Ig���;f�JLW��[4�+����#=�p�j^tۊ3�� ��D����/��`	v�W����;�Ş��x0)��4/��B�\�.�4��_�&@�-�p	�ػd4���m��u�C���5Dz��tŔ?T��g�[J���Z����[*��ؾkM+.}���_���$��[̆m�|~�H�(�B��{Thvx/��IQ�r�~��[[��-q��n:�$�N�Q7���6�� i�3�#��fȜD�S<��Νy)�:�<&��M���s���zgtV�V�2������U3G��cJ}�������b�fiB.�w�����_5��O�`* �!D��j%�4��1$�3��0#ѝ������*os���e�;��a$��6AԊ�:��w�bB�W��zlj����0tF�4�J��(V~k��-��T�_�]�'�ͦ��G�-OfIeDT���\L��k[)�����^~��.g>L��Q�ةaˌ�g)M6����\%dnH�9В��e�I���G!��	��(� ���Ou�{���l_��Z�_�S!C@��u����:�Ϲ>�r�
��-���O*)��.�ֽIO�i�p�q�$��˾���,�XsZx�Г"L|E�������à��y7��'o*�5s�Sf�V/�Fy�9q�t3��?��	�%�?}	�=�����z �����������gR᫅��eq���͍|/VĠy�:�3/ �cz>P��_�p_v-�L����|��o����Y6,-��&j�8+ve��B�i��#q�@�i��]?{ �a�[���e~E �u�(RW9I�Wʤa.�Ĉ�:O1�li$��&��(a���J�����ٖ�	m\�$��<$@f	Οm[&�;b�换j����B�/���ET����z��pB�|Y��� ���X�l��k����'��[�H�ou�>�,�ON���'�8,[֐��Dg�V6D4h����V�1�\K��q��g'坮����W��'�|\����|X�	o���j6V0ii��Bk�������Mc:�z�%jKm���2U�tt�%����3��[up7~����(�Т!�QY3Z@�S<C���;��.�\�s+ծ"��[�)m�:V͛#|˕Z�ˈ�D�@>a���n<���੧jv���-���O6nS+�#ф�׽ ���?���g�0��,|�.nc0V�)�~(��t�P����vpk:)��tIԞ;��C���yK��$�bI�%�������)����5���-"���g����9�`���v1}��'Sڅ�`�ؽAW���� �z?�.����o�� Q2<y��
���$��'QI�ŒL��w/�7�^���GsD=
-��p��o�3��>W��J�#�^5�s��A(��@PȆ�P���F}�ˏ��l%��v#����a� ��R �$����}�2��ccn�=��82����^mu��p(�w)Z\�;��ww+���Nq����;��������Z7Y'�I�ܙ={�3�K)A}N���?1��h)D���x��Ev��a�0��X3lΟ=߀�[�����Â6Zr%Ybv|�=v."os;6ːs��8.B�3~b،cT��n�τL6�H#�e�[���'«q#�|�NkSA�XE6��zl%=���b!3h"\C��{6�'�z�In$Z�%����zt�;��t��o߽8��y��*��䞷*!�X�ٱ�*�Koż'�����b���)�P�
ee!=[�1�8��-����z{{C(�^����M����ި�~��\�br�j�t�sN�-I��`�����e��x��ȓ/����OT9�z@D?w��|9f�}���km��p���L�,-����	��Q���]�N({�*^�����Ći��9l���v�P���6�n��m��Mz	�N���H�镅���#�-GV����
ѻ��1	����[�0V�� ͷ�]<�y�0S5���ɂ���?��0Lo�ݿ���,'�#��v�Z�������[��Yb���<�%gZ:��H9�bl0{k���K����j�iS�+��E1v�����]�q����L/Z9����4(�}���!O]�|��o�}�'�� jgԆO7�)Xک�l��i�?*{��9�6x���
��E�Ĺi!�r�-��??�nsB�.7�&�M�D�Fl2P>�p8��j;�V�Y�.YBkJp��.E�]���	ҏ�Ԡ�G�hUqGk�\yt�s�-�>v0f	�B��֖��ꆸy�u�.�r�,
;��:�$�}>F.��@� �c2Tc��S��Ni)9A���H��z_o(�:= r�|P؛?λ�jLpi�t�y�^NT���n7�T���M�K�e���M-�>P��9+6�P�?g���K��g'C��ٺ�F���o�$>2;r"W��W�k��	��݈`���`�L�y	�P�j?��T�9v�k�֏-\<�"��ڨ=L3_���y���[�!��SG${�"�ɯJ����v�#^5]��5���&D�U<����i�r;V`�s�
��{G���
����0����ބ��L�g����|�2Q�v�����}��_�炃=l��>Gw@��X᏶�C�{�݋p#��m��;fy0�>יw�&O\Rj:=�0ȷ�u�~ϱ��3�4�̕+{�t9�i'��)d�v�P���V���*��ظ�̔T������D�eP��F#7�]�>���Ǎ�Dԡ�ғӁ͘�����'}��2�r�2LG����j����1i�V�?"ѫ ���g^+��{3S�x�M:�S�ܡ�c���n�Nݖuۏ�(*cy�+:9h��{�d:��Yh�@�Z�f�Ew�$�^L�tԜ]�XX0h]���SL`mOB��Cr*#�hbӏ�-�w۾���nQ^�f���J�{1>+8��T��ZZ� ��Xs��c�{f����X��7�9U�cC����Z��Z��4�URq��eS!]4Z�y�eC|��R��� `�%�Ƹl��^Qg�m9����T��	&<�&��[�o��`���DfL�;MK>��n���g������V�bv�y������P;S�]�jED�p�z�&7�_X�6P�1�;U"4�[&-G���Ӯ㺰scN��{�YV�Hj�FP�;�+76��kw~C�^�ɍ�V3��p^� ͕3�?����i�O-���Wh]F~��[�@�<��^�zG3?����Z0#Fn�ܮE��<EJ�V2�bs<Q.���rV��f3�"�L���h��1C��)�oo�{�3:A-��z|��JutR�cpd9��7T������]�ϫČp[�`�Z�_޴�;��x�wϯ�=�WV��r��L�1t�Rg��3��	xd����^�\�E�CH"K�z��=Ҋ�DHI�����d3>Xә�PѨμ�yf�_�16~#F=V��/P��0�Y��Rjؑ��d�ӳm���y��ˤ����O��C��O�O�c%�3�o��iz�k/r؈x��%���SY��v��̔=��K���o���O8j�FN���fi�Rᩂ!6x�R�us��\��l����w�\d�4����UT[׭3s~҇n�ŗ\|�?�E�,9w��/�C��h.�����A����e�fb���$F��֌_�Ɋ�|41�+%�����::o	�K�����jB��_&)j@m�e�v\���x��_�@������0�y���g �J�b�lٙ�Qb��e|�bTО5���J�H�g������0�x�w�D��<?m�N�yЉ��ӄ0l����F�����1��5���=�@u'a��(.�*�x�6���_)q��͛�J��j���[���4pbBZ�����G� ���d���f�v���dN��\}�("b����Dq�4�`��7C)2H��Pغ�����'ע�ƕm�\�c�;p�%*S���?�:އ���ο�ij�㘈�������Dӻ�����`�Av^U�����y�Q�3���"P�k9�^vG��@37���E � |ئ��v<J�e!�F\�W�2  ���	P���h�U�u\]�v,d� 9����j�3�|����6��/w݆GK�������R���3�#(|W�6l�]�#Dm�C����L.&��>�q*�?� 't�}VRB1v�oɓQrѻ��>cyz�.�v�^Ptu2�F����~�����h�G����~�����L�^M��F���F)��8�? ����ظ�災#,��A|<П(���PV1@Jf����? ��@���ʘ�?���%6��]��48�������0���$�I9��)����vﲇ<Nd�C@�0`6��$&��y�[FQ�f�����c%;���ֈ���@�Q��a�=2O�k����%��N��OҠ�~f��%`U����w�i�_����{+�j嬎������܊CC"��'62�\Lv
�iSF�U<4q,}�?��'��B�`�Զ�ZO�/'?�@���j����hh�v��rh2<���N�e�z0ꓒ�nTn��s��~��G�t(k4��)S�R]����t?q<���o#U�b1I}u���u2��87��8`��1���S����+�,zv��`SZ�5����2��c	��B/d`4
��퐷�/^�H�0
�7��[�k��,Ab�`&��C�с�i	�=}$��n^���d�~��B��������*�����^���	4P�fI�D��}B����"j�Q�,�1�5�"b3�,���Ql��/P\4D"7ȼ��OT�������uǄ���I:�-���X.4t��L�7�*�g�j�Cq��f`A���(���@����*]+�����D2�O� ��$�a�ָ�R��@�"��#P���b�d� ��I�:�ݮG��ɱ��\;�ܹ�\_/��V��x�6ٕ��1Y�x�?��g�֜%BtF,�g"u��_�8g��q�(j��u��Qjd��-u���6��Z�R�#Ip!��(jE�ǃE
S��p�E�m�vb�\E�!� E6L.�����`��_�4���d��E/�Q��.�,�H�4�n��!&�|Swsc�yV����֎��k�&t��hi1dT(<;$zL���j�ͧoa���]��Mg==�����~V�M�W��"/�m��
V9��1�	w���4��9EP��C���ÑaC������k���a���%b���Z�
����������,�!��EaJ�_+���7?Z�{�S,>�}�^a�k�80��ml����O#�b�⿏��p���JI���o�@H�YHrr�_[��J�	#�����$�=�޿�)���>���gP�tЂ)N�����͟����l�������Et���� bӵ�mp$T9��{��)U�X�ʮ�`��g;�L�VA�Ҫ�Z�!	�Ղr���V����`1:�p"!n�
O1�aYmu&��f|HW)	2�d67��V�]`�U�Q�A��ڊG3!! ,Z���V���G��Ǯ�'j�����m�ڑ/=9;/���V���R�瞯8\Wk�P���>\.1k��Ng��f��a_W�J𳮢�p��Б�	���`��/Ɍ�\�&X�L(fA���%�����WNc&H�tC���i��!2���Z��r�Z��Y��=�l��.�\�+��-��$ґ��6�_��������b�R�;ʾ�^'������*b�#~��9��`����g}���V���HF9.d�����4}��[mgqtt�Q��?�9��ɼ/(赵����j���.��ʌ_�mİrZI�4�>��;����<_���@E[n�ڶc�m�
ϳ�f`��p�F��~�3[]�=m��[�d�"1c�;�t��l�����c0���������^����/Om;%]LC�j,�)O�����z����Ԣ�#m+�<}n�]e�ބLr@��Pf?��l�U|�<��1����P7�}c)��O���C�5ttI�na	�.����Yr3et5i9�o����'=:Nb�����s�3���'0��^F�^D�J&�E�{��K�6���[�OV�\�������P�Hez!��*Q��'�\���P_k����ls�o/Pb��͎j9�E�S��w�Ck���=����٣�C �iy��f	`�pP�p4FJ����lU�������7�g�r��L?��2g���������p��*)��R�)fAV��8��Fm���ݍę�t�ޚ���!�'rc��8�y�k��Yw`o�[8LC�)N�[���� �.j�]h��)�\���'p?�`��A����B�%y$�����g�����cT3ɒ��*��d�Òk�ˍ�1U��xl^�b��"M�r�Z���z)S];�$���}|��1�%��GY�XE*TH�I�I�z��N�w��I,y<�6�c�j��W�b� �*�x!�C0ʦ<��$�f�3�������z�xVC!��rЈ��0����$�;��͛$�50�ǋ6u	6��"K�l�梍 Z��f�^hF���\�{�݇���J�
W$�p�Fܿ�j�3�9�O�v
<h��5;�^l6�jG=�#�đ����~F�R�]�
���?�͓�(��w�yL(NY��{H�b0l�2�!�!��
Ж�]YAr�ǒ��(vG�s����}'���/Ex}�r�HTU���q^�{��[�"c���'�?P��;f�/�SY�_�����лv�t`�j�4ج9����+U%�,vȀwrd��Z
�~���h�H�>e+�� 7�t�h$�.!73�}����ľ�"��q�xí#1]�������Y���u�������۴j�C�!�~�������屇���r!�9�7YV2��p�M�T��/�"��yն��8�Efn�>E���2�1n��� �9Z��?��v��U������?�Yv����Ax��G�x?��.�6g�21,�bi�e�N��B��T��:٬���R%F*���9˝՘�G�d'A��dH,���dS�c�)�N��N�Jݮ�����B��?���6S�6R1�"t#I*u�<�a;5�,=�h��Ѝ���
>!u�z�Hȣ�2T��ڊ�p����]�\�}��\*���jSܴ��� բ��Jv�54�(��ڔ3�Z{03���8��	�~���#���N��V_��r�ӂv�� (@=�������n�{�a�|�$��t"8c��3"Dָ�-{8*��u�<�/2�(B0d	z+�y��Cn11��9�G���uؤ�f�Mˊq󐺀���о��L>�#u~g�5��'����m���:4��G��m0Y��k�_�_���<O���j��ck:� �9�fΝ ����]�!���0�~�l��u��m�&�
'F		hT���?=l�J�O	4p1D5�g�^�M,��m����łK9(����G�*X�!r���Z�zަ�c3X� px�� M���������G6���t�~/�Ux�빗�D�õ_<��c���}��*�f���o�����V�!d�:k���#=��b���⬽d��}qwG�?��q���z�=7�\s���pa>���yic��2���}o��k]����<M���E^G�$���l$_hp�?�äa!�x������`�M�,hm�=�G?\�	���|3{��A���i�#�0î�����q��Q)R1��HG�	F�g�k�]�oÚkٳ!J�F|LF2��l�Y����f���K�)?��v��	M�1V�;��7��XhYo�mP=�i�۬=hXC���$`
�(���	��~.0e�2S1h������";�Q_-�	�4T��}��b�\[$R0��H)�.kB��V�j�3�jeU�b��T�ɍ;��Pg�4mC�"�_��x=o��:k�"D(ɶ,/���Zѕ8JY�4W��\���� �6�����y��v*�����L�
 �r�k�������?�:Q�mL��w�R���HH�\��K�]��1o5&%[����D���~&V�������h�f��΃�i�йSn˄��g����}�e6�Y���ˁ����l���k��0�q�d�ď�:ÿ�t<Xz`螏�i���U'K�~�����ss���R�Q0�,�8�d�FҦ�����gw�Z}��Ai�٢SkQy6`��̻�8�ٻ&E$ɱ�[�q�V�!��q�� 4\�f�v+�@]���_�*�;��b��&�3I�rw�^8%��r*{��it9�o��0�����-m[M���w;�?g�Kψ���6B��BUZ��bd�	H��yc�s��*�?�.�}.�_^bT!��
�2���:^��s�Bl�r�� ¢>�\f�]�k���,���Y�&E5r�"������1��b��b��P���z\=�ծ>鳸�X���Uh]��f� ��qxx�b D�i�%�elDA�[��!�����!��i�|¤e�s�4f��XD\<^:	چL�B7�bd��֦m(H��ܙ���n�v����������vi��o��Pa/b�'�zI�s�B'w~.���t�o�,)/M!>���pIUS�יnv/3O�S4x��$����	I�ts��g�;o99]�*����۩��uIOCH��m�o�8rW3��-/N��D�L�~7��������l|S�ũ
s��]�7L���! � k���� ֵ����ID I���g�Q9�P��˿7X�;`�;G�{���O3�L�_��џ5��%���P=�[�rq�;��l�<OĜ�t!�Ћf��ٲ�S=�|5��qcA�Z`�KXD:í�1F0>T%���4똯�6�8�7��P�2M�����.FT�y|�����`3A�]M��KpX6b�6tC���u�dH���;K��9��������(x���M�����B"x=��I�Pl�;p��\ �L~�X���^�KΘŭ�%]��1g=�緍4r��rjѝ���g��9����E�GZ햁���L�� Ka!��Z��p:��ߍb)��������DG8���fg:˦"�>7��k���r�P���K	8f��{8\�^S���f�W�,�x�K˭P���H	�@5��9[q�]��%"��E�'w�V�X�o��D[w�nҨ��h�ݹ�LdzC�����Oj��|;�X���A�c��Dm�e�[�|�j�$�TCE�4�� �c�&�f�L�@��i]^G�{�C
�뿸�W<_J�#�dK�g�5/g��/b�&���VP* yC��;�l�HA`��S@1=�ՆL�e�gc7��v>��`{N[�a����jX��M�{�+�2�8�dg���-Q���)_�����W�zb�e��,�����:�r^�5���;�
C�?��ϰ$���4eQ'K���c�_�*��K�	�G!
�����ô��P	g�S�j������
�A���5E��B��;�L�7fH>1��؍�%O����˰���zSPg���&���ET/���p��E#�u�N����Q�&&P�I��)�O1^����V|䳡�e��muq�Уq��R�0��ʰ��+��ҥ�)`�]Ğj�bO���f�6�N~�f�u�`��ui�w�A�����A��m�6�CH@R:O|��_�Kk(M�k�ά�zRv!��pd��~`�~Sj�'C���Mq��Yj|�<��	��5��9 �m^Q\�LbwvGm�}m"�,_V�`��~�9�����rA���P���Y!HqM�L�.��b�g�j�P�:��L���NsV���:�R�}�Ψ�fe~n_����X��̣�z2����@s���	��k�N+��y�����M*(Z���tN��m�?��y�~1fd0H�^���^�Ikm9��1�=���1��g]��%��j�-�SY���ę0��,{��1W�3�C��
|E��s`����9=��~5��&����T��)�����v�L�r8�MB
�U��#�~���."�.��2��4����G�><�A'��p�����DC+R6�$p� i�~).���Y�'K��H�'V��v: �>�����u��@pr�.�T����&�Ўg�nA�qs}���u�,2��q�1it
Պ�ȥ�2�/jcq��hy�$~��9���@�G�J���K�������e��a��	8J!s���n����H�4���q���N��֑Y���y ����W�z	��n�W�l�������L���|GFU��{(�:P�I�]I�+z���c9�^�;h����|k*fx���6��r�0��Qb���B�;s>��������t��C�lE�P����UIZʣ^����#G���C�g��e���:��vb��a&��7�o�"�G�,,c��;���T0OZ������G[���۸�x�}Ӡ��g'TCD#D8�����9�l��/7�+�,'൚�Cy�r}xpi|e+I�_���MC��v�X<3cH*�;XA^̎�j���gr��D����s��L�鄗��D���k���C��~�97�qbN�W?DĒS67��5�w� ��0�uy!4T�/��b���� ����'kw"ˮw�����g�KF�.�E:áԹ�|��R����y0�T�ώ��4{y܁��zk�8<��󚸑�;"�}�a��U7ΜDLmD�]֟� b6�"'�W�+i�t���:��V�w��V���f��q�S���׺�O�"��6��;���:go�,���V�+��t#��~*����?���\�<n*MkE�	�{�k��d����vޗ׫���˵���q�@�W~Hu��1��)�hrR��VV �:3�e���Z�j�lvŧ�s��#�%o���U��}���S����+�N���Kt�)�?z�0��?�M��v�j���_���y~$����o�߂�}W�~�Q���N强�� �cy!��u�"m6�:�ԟ������`�4*2mD��3+��lo�qa�f��~��(�[��/k{��|a�R��y�c��"�
�rCw밫��Rh�d-�Ѧ����ve�h���~sb�l6�/�#,foÓ���<x���36��+��V��l���ҦbY�*�Z�>�R��!~MC����g�ԙ�uC5;V5h���𨿛���4u�ӽĄxLC?��4����g���c�rn��5����ݬ�]�7Ý!.��(J���T�vD�#�8�2�ݢW�,W�H!�|X��]�x?I).��������m����ڞ����J\�@;�_cT_��C��F��k��T�Bi��_	��wMX?�h�9��݁0)@��{�<vj?k�!|�4�IM��!�hȏ$�tB'�u�+X;
�(ӽ�����]��ܷ;!�2�l���6B�MO�L�P�ʬ�}�V9��g��r~:�S��PN��z��9m$�L��u���W��"V�D�w�:�����T���
�Bk/�L�ґ�ty�=�D�rBa�'��N��Z�j����J�C�d�?jH֜e{8Rv/�'V�U�A
�O{F��e�;Ĕyx>>x@!��ʁ��|Q�hO�� $F䟓
��]�t���IE�f�:�F���hr*�,qʑ{)O~�9�#O"z	X��Z��*�`݋Ta7�z+�͗��g{��җ�؋��КV!-��ҁp's��|���������C%Ae��wA�=�Bo:�z�Ɲ�}��K���b��^T�4���ٻzں��w�P6V���\��]�ñx)���;<blȵ><��<I�J���5-9;F��BC��o��:��7�uD�ۃ��x�D�5[�}�O�8�͗�E:v���\����a��3H;�|�rwU����-����C��M�Q�tKa���XM"��I���1�Wk�$Cۗ;��v�w56H˛yjۇn�}s8�Ϗ0����v����fw��z�N�zh�� 	X��x�M����*�̓�+T���(\c9w4�u/���dˏ0�P��'��p໌-���Fo�"���J��ց�s�A�s��}� ��-{��� b?���|�m "�1�A�}���U[ ��@�J�s�t���@�����3�Ƣ�D�B���r�2��l�P�"����6�2�p�'(�� -�rYK��r�y�ԑ&��j*ܕ6�Wo�]��6�@�����"c����óEp���>ވ��_�����9�X�4?�äg�GAA졁��&��jQ?$��1�D����ו�9�]؇�WN�I0�{{,d�ؘ�/�x���V���ը��7w?`Q|�@�m<�p�,�nOX�%�s=��b�"�aY����B�KO\%q ��oqU>��+����d���X������Z�v�H`�-��):�3����,Z�Er�r�$);]Rn���4��3�������u�tF�uwJ+�i�q�mD�jܯ��_�����NQ��&.C��h����p���O��%����˵��U�E2���VOs������}���N�2d3�����A����/|�.��y����N|;�+�ȳ�Z��!R���/��E����JaN����x�fg&��cK����ܛ<��.��tƪ=ļ������S�M�b��Qs>X�|��T�`a�_��k���7�����1X�����{)�1����h0#���f#�����]>���L��Ͳ��(����^w���7Oy�~�Fd�i����x/-� 6�8e``R�#<��-{ܡC}j����E8�  QX�+% u4��徵��� Ş��Fy�ss���8��q�����^YO d�Ӂ6WQ�xP�.�]~A�v��N;.
��~�m�y�iک|�v�rE�L$�Uv8B.�� Jn*�c�g��V��<�	o���%כ��wOȏbh�ǹ�F.jc�ݻ���;V��g�;�������]�_�J����GF���c�g[H��D��M��";I:1]7Mu�L�s� $bFZv[�����+`��d(������;-�S�"��@�I�QƖG�#ʋ1J�`!�T��Ґ�˒�-�˓@u���$��L���7�E��iU�f������*=�e޽_���Ȼ�\��@!���I6b�2���f5�8G�� 'I�p�1i��C�%Ռ��s�������v"��,և�D?�D�R��;��a�$��@��� 8�/���T�c'9w
����p1K(��j�ʅC�"�M�j��o��i����s���m%A���1�Q)��9��$���L]��dX��3)�������4t�BO?���[M��я�����S��m�;c��!-�MH\S�&��`�φ1���7���jh�o���Y�˹����G��<����^W$�AQ������S-zF���.�w�ԖG�a������,Lc�4��S2��gF3��WyT��J9��;���&T�6���� �c�`��;�03��k�����ړ��*��a�7�s�Į�|�wc��J�t}������ʈL�x5z1�_I�v�������SI�1+�o9�Jb�;*�l��T�9j�Z\wr�$9��v��u&��գ�t9�K	�;�; �c��`.�H���:L|� ��`:�Z��<���7hhRc��\�5�^�
���(Y����X�d ��>�����(|U�RD���ɬ\��)�ޗ���z�b��X��1C�p�B��x��ĭk(��<�����<63$��_��D2zTy
J]�[��^�)���ZUؖM�x1���#=�H	J��9�XD6���f͓!�s�m�#����a�G)�����14����o2��-{�i�acVc��}��	��X��Ea�a
��&�XNR=#S�o�[>�*��amxg��//���^>8D��~5µ.G��1u���t�����j�hj��#���M�X�[꛱HFnn0g���P�:�a��0��7z���X!݁-?��%���'ȷ�|,p�+��lhz��8�+̥���oP7�=[���+_F�2����8l��l4�Ud�ٓ��~�-�1������aq4oq�!oEm���_���I�(�/1��⨛�0�	�G�7���Dv4N��YL(�v�9��4!_�� ������`y4�/%c���r͇hR
��pDT찪)��k�e����4���>M�#��`v���0fh�Z�&��l�)�0��qp2A��X�#��u�k:/��Ze�Sa�9��;�m��������~�>�杋����p�$(HsX=Ey�����%�@C�
b���̖_[�B[7����'>(}0J�t���l���0̄�"�й�6D䩔m�F�j4Β��HvuZ������I+�4�7�^]��A�'##5�7O�M�T]_�d3��6����#8�h�Lou�NE(O��Ɨ�0M���3W�S�,��C#=C}5�ȇg�8��R��9�rC?���KE�V���2����w.�>3�g���#�X�E~jnJ��r�|��.e����b��n��_4�<Y%��۵���\a:�e����؎��_�M�Ϟ#��o,���G�z�(�� r���	��
������?���
,���@VZX~[����T��=�;�kl5^A����.�0����vR���z��:���,�Hx����']̜�oyK/e6�	Ke(�:҃#�i�ҲZr&�d52Y�7%����[ǽ�N��_�-H���!OH�����x����C=4
^�\��UN��q\Q�9�9�iJqG
�M�_s�=�>�^���_�z(n���d=\�0���1�Q8�쀢�f�A(�aLU��,L���<H��ۖ@�+��P��J��� >��BAr�VhL���Q$BCk��c���XD���yA}�î���oݥ����i 1	�����`p��/W�LH�a�vϟ`�}UoS�4N�-�å�>���W�ݴ���H�B�=���"�Zr��G���y�&+��q����m�GylG=����%J,����fG�v����>�&O�_X�D̈́�eS��8]/���0�tSk4u^-`���&	�\G��Fہ:�b򨡘@�>8P����g��"4'��U4Q�AO�CR1���>I�|�_T�w����Km�*3��GI6�0\՗�Un�����ٔhՎi���y|?]ws�6K�|���k?.]�g��0rع	���'����z��osq��bl!��������_P��K�r���s�x�N�o�r�݂I��N�<l��S.�fΣ�܅�S�knWI��op���&�A��{ԁo����s��#=;%�:���C�<��6�h�b+}�Jz���
Kо�Z�V`��10���>�w����
;���$�s+�:����i|G&�W��V��D��}?-;!FW0m�|SC���Y|�Y�n���8"���f7��/'�^� ���ص�P�mnME�}P��XWK����\�ʄ�oj(EUc����m83��m��ah�m�������@�`(K��L�L���x{��e{�b�ך(|�p�N���͈ɧ�B��~ȴ7���oS�s��{œ�̳�$YO]5��Ŗ-�[�Z�q�d��;���(�}���|^�@��q�A���@w6�9����#Ux@� ������������g����Y۲�̸���:c�UM��²yy����(�~հ�����e�^����
���èp�KLqk�n��j��w+�1������c��˅v�S�Skm�B�)�Ђ�#qf��i�55�ѵ�����&Y���U&�z|�7g�4��H�#�!}}<.S��v�h]��Hǖ���Wb]]� ��p��I�g�F�n�Gž\�oT�!�+�g��܍"_�%����2��țF�_,�1Gr�<�}��xk�X�K���~�r(�d�	�{Y�ho��G|fN���Z)�Ǧ�#de9�\��	;>���f`S����EL��U?�S��B�7��e��p��~w������SU,C�_�]v���jw�!��D���m�9X��i�@H�WH��~�����m|ʍd�~s�#������כN��><"/ �m�'��D�$���\� �?G��̙es5;�b�~3���|}���Q�l~'o��|�����08*)�Y�%��@�߷9��{ŉ�%V��ƴ��4����i%��;�y�N/���:�8.^����Q���f8�� 4d9���I����.{��5����
\v�y�������,M@�=]��f���hy�ԦպF5�����;����uH����I���:bQQ�9N�����ß��|�Zo����հ��k��וu>���ǟ�h%d]ٌ��5��v�	�u�i`�oU���|8�,���v��|ђ��\�4�LUA ��1z�r���!�g�Q�I�6��I<]�����[�.�9ʪ[�����M�f�yÕ��q"�Q(2�F�	�����˻2���·���+��bv�|���X�o��a&����x��k,g��d,#�K21��A,���w�Y�J�l�PP������JHj��-f�q���0?�6i�'Q0���
�%e���Y��f�~��w�c���;�!e��3@l$�r��׊H�ټ;�x8��(��6����Q���Z�Sl��X���ؑ���;�����!��Tj��]c[���4�+�ޒ��d��b�Kz^�ļ�=^�#���qh��n�Cm��c�r�E3�<s^�9&^	R���UKo(�1�D	�����z�b�dI�$��j�����>��E��@�"�4س��r�X��5˺�N���3��b�����n�v�1#c�^x����r��
�T�����OP_>^Y���T?M�EAt��{F���֧(�~�+�� ��Lp�V�!
)�t��/[Yo������(G��8O�1��Vd�1���	4��! ��w�tz�t��cqB��5�aZ*�jU drBi8JZ*<�f�QԮ���;{0zSQ�1q_�%S6��ׂ!'����ȥ�P�q��۾֡���?E�i_��x�Y3����e��u�_.�>�(B��D�&�X�Aj/��$������TTĊ�|�EM�W����/	��,%�'Y�T��?�i%�P�}C-�y�8��[ֵNW�+d����٤�#Y,ꑭ>���2Fd2c��YݟF|����L:*.��b ��3 ��i!��S0�!��'y�Y�*!�ɑ$Pk����,�]��������|�T���? J��NH��E�5��E��.�>��Ɓ����l�a��Oh�a ��ȕ]�ќ��>M� J#}dÁ�T�00XE&@'��L�V�X ��P������X���d��:�O$�4��&�0@|����r����x'u�ǿc�dM�yZ6�z���fZ1�CI@�R��=I-T#*�$3>��
�9(a!��	uZr	�ʨ˱Fd!� <=DQL���c��>/�Ke<�)�X��-�_9�Mit�a�PkSjjLh�)r�K�uW��
F��R�[��9�G�ɝ_ğp�)(����\������Nw"�����Qfrg��7d�y��:�S�nt�� �=�V�<]���b��x��2�-�)��Zp^��J)�D��<�8UT����H�+�p�"JC>�Uy���A�,���b��PX�f�D���:�h��ݎ%�S���eG��jUQ�5KŎ�KV� ��gv3�K>T1E4g��ZF�磙~gME��h�$&n",����֤�7��ݙ����3�yz?��'���g�)�X ���r��ꆪ���*.���琐L5��kƪ-��:l�b/%�l���#Ʒ�P�N�[�*ʏ��@��Z���h�-�x�)7� �"2����V�L��/P�~+7���a����i��Ԇ@�����4��JE��N�.��g�|r^��g��î[i��'J�s�<�p�~��*2O�F���~aΜ�g�Θt��@����jrs��j���F����8�,"� �?���-�&p�"444 `�B���\W�]�dB�=L����*È˔Ýd��!	G���)�����G�;8G��[�Nl�۞L�L<�m��$۶mۚض1�3�w��'�ԩT��;��׷����^)z�d7�Zt�M��K�7$8���\B��������WF�%N�DS� �W��gˉG��k�fz׷�#"��dz�d�`X�������wM�ݑ8C���v�6R��-�=Z�w�jڻC˄��!q��@҅2����5�a,e��f	���G�z�oˍ@��"�����#���Ju�A}�9>..�ޞ��'Z8A�Z��tx���G��<��d:[�/u+�nԉ=����Jiee�d�8x���_��$�P���0�mb�!y�9A!�/�S�t�
���
�^$M�r�a��00 B|�k177���H
�%nh*L�v���T��dtl����RmtrS!@X�б!�;" ȑ�bM�(.-M�׸'	��K�L�K}�Av0�$��G"'���UW���LA%��eg�{�`G��-�����u��BW������?�Ч�4xRcLW��w�[|cD����B��y�� ���a �T���D�A11�_�Ӑ`� BHJ&����,T�S����НVſGW�2����s�ϯ�0��:`�)��j���)��Z�Nz0(L0��7�熌."4���p?&�>�,���O�x@���O�C����as)I��7��Ȟ��`�K�qN],VM�!���N���DC۪ʈ��$(H{OJ|�+fۦ���o�����5����q�˙���W[wnM��It�Mny�r�U���AVS�"(�<+�ᜃ�t<�����]�xu��������锭���s�p�"nw�D@�nS��SL���i P�3��M%:p�\7TAE;��jR#���CRwx?-dp���Zz̏&0�4t��o�r6���}<O�j��
���7������}j�NM����'b �YDpz��eӝ�����#��I+���;Pv�'�e��󖢥�~���Dڵ��41M!+Ɋ�?���5�i>����J�@�1n�������s7�|A��O�A� �O�P�-�k]%r_�ȿ�}@�<��k�p�>����rk&�ҹ��ܸ=:愶y��9�QL�-�,���s�(a�J�#뽆2ಀS(?႔��9�"Y�h!5���$��E����h�y��6���H$�(P���s�2��y���Xn���c:�y&F}�)kJ+�r����-})۾�O�,��2I�JbP�\]��(j'�pJ�̂������e�P���w΁���,rU׭�rx���M�,��AO��$�
�X����A������z�;���8c�g��-w6�(��f2�+��עc�3ݞ<;2�J��c�����)�K�ժ^�S����|m4�y��	�������/jZ�%A�bnU��	nJ����Rڽ׺����ng�O��/-���o�N�]	�'���Jܓ�^M"MD���	�ь[E�I���<v`�o��f3ny�9���3/���Sc�BfM���1N���4����ު͇��{��5<=�5ng�;0��{��/ 8O��v���?r���r}�����AwȦ �)�����`���=�ʛ���'̝1��J;�������:yH�ߙ��r�s���,��؛��ճ�$�σ  ��'�_D��G��@TQ'\�ϊj5�V�8����?��e$R�7^2n񻽵�U����[3RK[cI������կ�<�.��������5�7g*{ktj*?��h6��S�#_���9�� ˡ��;��D��~�"��JW�G�����KR�Q�z��+E:[d��E������,��)��tٰ��ӏΆ�d�~�8Tf)��uxh��I�k�q��4֩?N�c6��^\Y�u��]$)���K@5d)m�X�C+#4�R��[`�T�����0���H��g�S�!����r�ѶORc�U�ժfG�RLm�����uآy��T���BqdP� 4b	Ԧ_1A�:��$9�燀��L�y�;o��[o�Ȱ_��r�a�^9	���NKq�&�0��$��NmT�����5=�����M��y��X���r�saJ�
k5yM%���d!��5���`�8Z�.3��ǄS���H�P��c1��݌H ��nM���0�ڽ_.����[��W VȞ5�?ʜ���/�#zp��"Ew��&�cE���'�PI��4����?6�n��
��a	�"Ǹ(���="���H�{-�C���B����)�YO�j�-��7$�B#�(Q,8HF8�D�F8�`��R��	υ� �#3���:�q5�$�j�ҽ��a��tx�n��{�<^���QJ�@kw�'X����p@�P�3=2Q�O(Ø�0$p����������Z.�6M;��k��o���#; ä�C�^�ls;K%d����x��l�y�-�Fu�
�寴-�T/k{G�U��«̅n�z��-��m���L&!�Hǭ!'(U��)bte�#��H`�g�	ոi�����N/��(H��grњ�A��X��"�B�� ry=j�I�互�}ۢ�?@k��u	QBw�[i�z�;?UDA��N��N�l�{~�9�k������:>Z�6��I��
���`p,��N�ǻ�+����rWv�1��O��(�������3Ո_�u�I0+M��~�+B������~�R�y=� a5<*t<��D#*�S���N�;�4^�����D���&'�3��rN'�B�m�@�v-��rPz���0�(r(w�Ǿ�E*��W���3&~�Ab�[i��V���ѿd�m��a�b�I�a�J�.�Pi�^������m� ��s�t6WC:�3�!�m^G��lx���.�J�[WO���0�ѥT`(�d�#�q�q|���R�� ﻞӾ�{B��z��f�q�yY�M'6'�«~!7�&��ϔ�tCȒm���k�E��ԕ��#�0Ps�W���bbx>�V=��=�n=����&Uz}���5�=tc壼�wC~}��Q�ߤ~7���>�4ːW�7W ��E� *������q6��)A��A*���]�RV��~�JA�C'�9ߞ���rșW��U;��*T�cԀ�b���Gĝǐ�����:�fWo�N�HK-y���MMd�q*�忞>���1����w�pq�[%̞���#�_�����2ZX�>\
�w�J�3O�����)F�ۡ�UT3���<��Rf����"p��RT�0�+Lǭ�3����od�P�i��Jwp��"ֻ�@��N79�ņ,e����~��)J������v�xY:�&�-AFP|��F0gR4��$�ȓP��?YL鸪��h��8���e-��7�h씵\&�j�:k�*>��l�T����C\���B#�F�!6ϩ0Jh>N3��6� �H��nO[��6Cڶ8�F�JL[>���;ο�h+�0D�g��`�����@^�3�͞s��**���_�h��=ϡ ��4M}�� �s���a��LE���DNZy/�A��+~t^*f�ʇ4��T��.�OˎY�������,��(�E�g[C���4i�hl.�M����5O�����I��8��PJEwx=�gz�k�@�UF}T��Y�Ш(�� ��r�U�bJ//~:M�^�*Uؓ>���r��FZD�}K����9wmT2RnK�Ȝǯ� �_�l����ƣ���/2.��!����
y�2�V\�m�	[�'{�� �v�*Zl�?�����oq�K�|S)YY�ۣ뛛�Ώg��؉"N�)\5�)���b��]��~�{��?6��\RbC����
2ѯܰr�������ch�U�b�+u��8>�ө�� ��e��y�7�k%���s���)
&�@gp�ٮf~ُ��׍��xf?�<���.$���O\���b���ܑ�����)����{�T���yhS���yݢ��[O�S�5"�<y����딁ɜ�.#��Va����֪��
f�`}\���#���	L_�hEhŵOZ:T�7n�'�F�]��S��ElO�B. ��JO8����8Ӻ��z�a�����Ew̓v��ِ��*�z���~Ҥ�޲!Ve(����q����.=2&���\�E)C��j~A�Wւ_u����N��g�W:|	Gr���%\�j�x��s>s��`H�����<Ʈ�6�X��Kz.�	.S���&��KwҪ��kk��<��u�t�����HLy�����YN��]�d�+qԅ�-�G)Ygۓ����q�X[����G4�Ap1���w��B��O$f�9�-6Z��Q����S���1GV!>�!~w�POĦ�����������+�|mp�f��/�@��)�*�'�����$����Ĉj5�ua�q��/�,�Y�����\l��:�/ PU�j��E|c�bHK������&����㙞��T�D�j�)*��Z��^���gO#�t�7A؛:
�|��F|Ԁ�Ä��C��@)F�n>�ڄ����>����t!��Qw����TԖug�����X����A\�I"�w�tx��D��]V���
�4�1߲��7��h�5kt�o1�@��i��^�����K�\�u9qq�;}eFզ���*�b�6ł�I�i̢(�Cre�`H���pjۜ �@��qe��Q�`i^3�!�V$wS���V���{U�y�� �Zv�<�Y��"h& ض��\��|�{}ɼ3�%���avP���P3H0�Sj�A:�Y�Ȗ�{;ׄ�gO-tO��Nv �ݡ{����_� LϏ-\��XGX�N�"}��t��t�
j�X#�!7�a��o�5J�+���]�۰��:!{}��ۿ��k��vٷZ�-�����>��y��y��w|-�b&.Ī�8�٨�"	�H����b �l$,�G�
>��7ՍF��m���Ȱm�h�_]�_��Pud8h@�~��~T�7�e]�dltHQi��2Z� a�lU�1�<UV9Ȁ�^^�c��wB}/��,�~D�.�$�Za7sR^��uםJ'�cӾ��5`@�:��[�����[�6�x�����|P�& �[W8A=�e�	zz�jX�*~��HJ�
�ozȱQG	�G�X�Q����H��}#�ဖx�ʸ��Z�P�u"
,z\���y�>����mx��\��o6����z4#��ޓ�*a4M�s�xr#���Ø�{yu�"���CL�(��˫��LE�We���ؖ����39�֖�3u�s�YWo��g�j8���P?���׶|�M��c-9���Q��f��e>�?-�#����93�}LNJ���4tT"�����%��x;��M���;lh%t��%b��s���\���=���;2��Î�ﰣ��=�(�	��7���Ǫ�!:���Qs���YY�Es)W�毷���k�
D0��� N�����hk�ʇc��ks�>�� �Xy����`����]�؈�KƗ	����Z����==.�h��`�H M۫h3NK&�O�hOP�X�T�ގ����jM�׍U8_� zA,8Z8˷���}�RA��c���,�s�}�oi���W��-��e|��d�cmפ��]X�i�w
�.�M������e���I�:r�=nx0�w��[���aA"�|_2���v���;Q��O1 MЈYp�?��zA�"T�/�Dbx0��F$**�"V#�D�=LI�I�3N�XC	��@D	yE&�����#�πC��[iy��L;QG��)a��F �v՗�(@�XV�0JI�)�uM ��FB� �E������lЪ����`X�ӗPJ�D[?(o�;:�3L�7���9�O�0
�]C�1���Ֆ=}�	��ӫ��^��R�{��L�t�؂�)�E��k�iH� Y�Ux�
F3$j��u9@Rk2���ޓ��G�%���,)�Ë�S����,���Kie�8��v��Ap�)X���f��d�0��@����N>	�<]?�``��B�ŉᴣ��ܓ{�2K^��m������q��謝B�����L܈�ⶆa�P��߁xo�n^��6��<^���K|���}�݁W?���3�:�TH"8߆h�J�Wy�Tw��[\�?�e��@�w�%]�Tdq��'�QG��i*��ǔ��A�8�QDR���C�n�n�@Cdy�vݸ�%$$�g�\�ʛ�P���<=3�	D<(e���/9���<�(V��}�D2����L��rL���������(��S��2�GX��p2�b�셇�E7�/r��c�Y�f��GI��!L[��o�k�)r��z>�:�/4Y�wuc1��mp(4g�"��W��r.�P��/�M�l�2D��ֿ��EE~�A�+Lc���7��4{��[j����U��84���17�������y���l�l+ڟ`�����
����)"��,���O'��ε�PRo�]��@/W���թ�����?�vq�����sf2�琣�ۄ�v ��@����,�~Y{)���)��C����g6�J�qY�	P�Ы���r����lo�2�ϛ��,Qt�tA{�6����`���彤|@���|��ha���!�AK��h:x��$��$�!q�G����U˙��Մ��2�	�3��f3�K�z`�#;P���dmփ��qڗ�f�����aQ]���c�:���S�k]^�졟��M��P����D�[�B
��b��VY?����a..��-���ׇl�A?�A����0l�A<��2�t�6�}v���3-M�-O�H���.H�ޏ��ʫ��L�'�`B����	�$H�/k�|�k��`�XdJ�VKgL׍
85�����"�Qp����n!zkVV
��j��PО��k/��غ�ۺ�oۺ�2��1&벦������AA�� #<�\�
�b���!� �Q^��yP�f�g�_� �lE6����5�N" �3�o`�E˯"�/§s[?�8�)O��2Dã;ER�Y���R�'��Ƕ��N�R4����Eט8�1�k�3T�'����=���ꀈ���ZZb�kRAX�V���~%���$Mml����`l^lDA��Ht��!���	��͎�0��a�_����+���L=�-m�*��pÙwE�������0>v"����-�U=� ���j�5�ga!�s��)�($�u�z�i��0�����ˡ>=�*}k,��:0��V��d�H?,ʳ�MZ��� ��Y�pUm��:27+V{��w�����.����@/��~�Z�@%�Aѻ KRc�cW�w�ͬh�:�l�Ze(���+x�E�<�&M�8Ɔ���gp�7��y���� �ث���i���3�?׀Wؚ^q�9<y�<M���,�k?���te�7i(�AԲ퀛D){fs�_!��t�+��W���g5��
�=� ocQ!��N�~E�8my:k�Q<>�8������^]�[U��HI��v�ޣ=!c��	k�*-��^���<�:-�KDhg��G�L�|X��R�YB�x��2�#1�L.��E�Oa:�]� B*ߪ���]���h1���U�S� �t�5�`©�:���mEl ��ɫ00{�J�Ʀ��8�)G½k�(y�?����lgr٢�j ��w6;��{�4�L����!iŦ�h��EB@e��x�粷�c�5����5�xY�ph���~�awN�Vy���F���6�H#s�)�!-��(�cւ�O&�eۃ�e�B󭨉�4n#%UUO��`��E�ā�3�u@ �1��p4�U��^S�!ihp���r��;������cҼ���/{v��$]�:�H5��p������Zt�&$힤u�φ�`k�����%��+g��)��v�-R^P�*�����K���;�g�F���<��h�v���[���f�|P�M$�Q����|��@(�0����6�m�>���{�q7��И8Q�Y
.�o���R ��h�Bĵ���st��|�Qb��?��ߘ�{�.hX�=�����(.���::��k�s����[�fE1z���^>�v9=��RQ��/���8g�|��t
���b��@�x�n�����9w�]LY��^�5�iw���*��,���m���q-�RVȖN�W
��3��C�<�/`f\�-C)��qwy�B��Seg��)��q&��Pd���3�S�Em^˚Z��a��8ˌT+z�ĵ�
�h�웠�fod�}�e%�MC��zXմ�����3���֢v#�x^��D�L'�ܼL�-M�n��e{��`he�d���W��'}�����)���V�廤�p-�cy�AZ�*�@�ig���r��y���ǟx�2p���zjq{�/B_�`^�G��!�����AF��a�+�VM����lbx{KRl;���K1+��.�8��6L2��o))ю!���z���Ao>;��\L�X.v�nF=`��"a��X�E���������]xї[ލ8��_sB�K�������Y��̵��U}����D�ƞq0oU���T*�,T��h���,K�z��0�Fw�x��򸾑�qލ2�G�G#��Z�u�r��M�Q�"ybuT[D���x}��5)��I��,vt`�s����'�}��H!�~�&�AƔ���,a`�r��k�1��O��4��.����i�E"]<`������ke�#�X����iZ�����ܠC�\�=j�g��g��.���{�JO�c%��~��%`hԾ7aL���ep�����y7(�
��`'�m�`g��=YF҃Z4(C!�+�g�����/���NC_�d�Y�X<q0��ԵY{����%�h�H�qɿ�K��d7������ś�x>�_p����6�%�qy��=��RQ���Л0�|%�������ƛ�}�/�-;�	E��P}���3ѕ�������u],�>���?GV��_�?�Q���B����n�\�z�%�Z{Z�=��v��^���;���"�W=�&p�\csR'Uy�װy��y[�<7�=tJ#�t���ɍ8��Yq�K�D�(:7�~g��JD��fپ'�,V��|qdG{���[y;Vc��Ʃ��}����U@�76=ӟ�g�#V!�dw�y�����D��kI`le8�u!a����������GZ��R��-��N�՛���"u3<3{�<��QT�Ѭ�.��0
��I^�K%����K+�I��O��� a}��U�1�-�G��E�l1'AW�ʪD8�<�όe�Z��i��,k%��5��=�&���cCќ3���Y�m����ug1�Kw�ԓ\n����#����m�ࡧߔ�A�� fo?	�o�`��>�-ZHru��D��ޫ��J]o�B�T�80|N5�?�	�7��Ej��|�-����&X�a�>�>��ML�@8�,���]�I��ke��K�ȡ�����Au5�4�U1}�Z�z�#;zpB;� ���0�����Kt35�l�����^͚��D�>w�
���3���v͹NсQ	��wF�P#�w)	�?=���o�%x��z����:oYh��6�֛�c
qE5��U�`���2��y��`s��}�E9�~' ]oo�
�֒o��/O����RrʛI|�tXRBҁ���Å	�vhx~L)��[���߾�G:{,�]�.$_�$5xk꜏�q�N���*b�3��I�O�j����R~W��N�E_����@��c�^�ZFϲmS:��5�*�2|.��W�@pL͂q�H�_ݞ�X�"՚����g�1��Yį��F�����ґ⤎X"�;ԗB9Nq��T:��ј�5�r6�J� ��mW�VΝ��V_~���a1� j�
�� Ӟ�G���D��d���<L��'��F^�K	�;s�a�%�  %�vc;�{y
A��a�,�-�K�tZ~bQ�H�"s]yu�Ԫ筂&7��ɻ
ѽ����"�/�f&P:T����]�I-�.��y�P"���t���B\n���#0Y�F3��Ct�϶�AD�{dM���"h&��48�Q�q��s�,b �3OOI_�NK�m�·T����z����mw�2c���	�;�%���s�9�Z $4�+Xg��D94�9�RM4(�Л_��?��3U~�x���J�밅����eb�4�dʀ����;�	�yD����U��(#7��[�(��f؛���
N���9�ԁz�?k��Eބ0U��]H12\�⣔��vf��X���K)�.:͏�7�ka_ӊ#>'G�a�Iǭ`�|n0y;oH��j��"��㎯��v,a���]��N�mc�}� �#W�.���
P���S*��ùD��ũ����rdQx�^�_)s�@��9��:�?�*y9���,�Y'囡��ņL+�ni��k?���O0��9�y�?�^�@q�b&9��4z|ϻ�GW|X����h�^_��7���r�k. �TJ����ke�af�y�̊���ti�,&1���<��Ac�����5��v��o�N�v�WkQ���u�m����*-�ɬUD�˝��`��款C����Q���[.�������rh�Lt�-��w�� 9��dTR�!��%A+�Cڗ]Vْ�B$�fށ��M��)�V+�ua���{��5>N#�Bqee�&��ZH��~Źa�П@��[���
�3�.��xe��;����wwo��)D����8B���{Z��N?:3�h�x3��pn�rC{�TZ
��Fy̍��RD�ϱ�6^�����
hX���P_�,V؝��'���Ʀ�����j$�3;�q���]bȊy]d�\Y��+���n��hq������-�E��c�Bͧd��飼�H�Ƅ&zo�� To��"�g�L,��X�)�Բ
h�gn`H�y��<����GR@։0���+�"î"��P��I
�X��܋�=��0����9%z���y�m���k5Н?�23RG�V`�9,�?�L2/U\����49`f+��ׂ[����tQm��:�J1�9⵪o�S��߲�:���b�AT���ɟ�%w;94�K�"�?EM��q�����4�����6tmx�Mt������2= `�� P�jX^ڈZ* 3k���TDd 5Ԯ��t�S��'v	�ei�|���������VNQ�n@�n���^��=���զ�Ǎ5o��ea�&G��!s���J|����{��)�F�8 (��,�/�?eWhl��ZE8/�v����I�r�}%]o>#((\�*#˪V&{\z��T���%N��Ö���ڱXp� kW|jI�\�0T!���R]���t3`��		C�y�����K�2�A���%7�[��	��ӫ6���;�&Ƴ�& �="(PZ+���\�-���5;nZl�#� ���ٯ2�:��A\9`��5�<�Rjꬻ'�Z+�o�������S>~�K�Pkפ�K���/���q���tހXk� +t�����BSE%�r�[�嵺�S��\��C|�K<�Q��E6�lGT���4N@�SJF.�?�5��<��|j�W#Б��sd�x��r7�)�To	�h��+�'U����ipf�oң:@k.�<��[���F�˙'g��J��{ ��a�\8)/��j�l���-��Kd44�]�	~�e}���gKf��.> >D�t��Wv-;�	�y����B��8����U{#6]����/"}\�f�}��hR��(�̚�w0ye�\�^K�o��-Nk�z�P��F��K'΅��dJ���|@`���V`�&[�
Rw7s��7r��vP��dĺ�Kwa�V��� F:[N���5(��2r��;���fhAa��#�~De�n�?���;
����fU��;@��>I��9�3c"?u��{J�w3rV��+m��)F�i�\�U�@`��MZ�$�l��2X[�-��E�V���⡁/q�ki2 �1�����P_<z\%��<[����
����v��!�h�t�ܐd���S܎`�$Svtkqp�L���e����&�4�1�|ֈ-�v3�db�71;����\ǒHp�zw�3(8�$��Аa���c�B_�w�A�$(���,��׶�hf���})r8�3���f�hu}�~�G7� �7[&^�04�ÆLZP�鄗�[+�Q�G��]?��"�}��u�0L���9�c�{gc�>���3�?�)0�(1u3�� �wsm�7��Z�wb()UA��VNsΈ]��tq�_�g(��j��{x��t�!�WY8�.��G;�����z��|9vo?�p��Fv88ӴFq(��oNNl�*^]��"��޿��nv��"��E��SSm5|"��ĦvT=bv�<���L�i��!1�E����(��]���r�nno�,�Q���g=|�fϧ�؏�U�5�\��0|A׷���YY� ���xVZ�!�@3��;� e�3�ص���Ъc��z�#gi|?O�x��^)�%!6�gO�G�"�n��V�gX��
u�.�v)W�7O�-}�΁ZA?9V����J��rfΩ���B�wqU�?n��F�5jp�it�"y
�fO|�m�R
�Խ�=��������8�Sӕ�0|�er��ዋ��H�u�iJ�X�I���5L-��c�d`�3�2e��^^S�2#�c #n)��"�|�xu��gz{;1�uZ��X��ҭ<_\���)g�D�����@��ո_�)>TA�|��`��L�i+��o�҅����8Xgc�K0��B���컷M�����]��Z��7��Ƙ/�����2$�{B>���ϔ�Бx��/�"���3r��?*�_��Z��e�Eř��� �G����*[�'T������_h�A=�h����������3s
�7�Ӷ�� �\�!4_F��J 	&(6)���K�Ǐ��ْ�Q(F�5᭼�si���g����c����۸�+�'ʗ��^�NpAs�Y�:��Z#E�2m`g3���z��	���P��dMbWCIP�2��Sd�HB���rFnlh�N��]'_��w�טh� ���ݸ�D�B�=�P����\D�E.���`q�2�跴��M�AM�Tp���5�������%�ʪ��C٥#br椊UB� ��a�7/��y9ό�c�zp@Pm�b�/���oT@�ș��55tj[e����%q1V�&�՜���(�����k�rl��}�VٟaAQY>���` �4щʹ��Qr�?���Q\N[¾�(V�� ��,:�o#.�-}bǦ,��,����w-�X��@�t|�E�Y+����]ʬ6�n�w�`={
���R� !��8�'{�����U2\�Bcf��x����������#Q�N �i'�?���ܪT$�	cM��#��h�7f��$8H�B6���\�.������ɒ׽iD���ϯ��Ӊ荃�V��@6d'��v*&��,%��6�9�U%3��*�J5��eȚ�x��[�z�gz;��(��#ܥP�b��C����7��?���q5o(ʹ_����-�V�_X�Q�p�}J������v@�?x����{|���˷wE�S���3S��b�U9�̓Y�P�^Ʀ�&�
�s��n��P�Ow�~1��g2��Z9����,��M�X؞ϚSz�<�Gu%��z��!OMG%r�O*�����;���tߤ����չ���Pu,�����nݡ��r���̈�����2�p(� hP�o��Z�6��r���\bcB���_W�g<��N�3w�ji���{t����Qt��GEv��aVI��1����v�6#�����Y��>�9����ڏP�?��z~{{���������3��������I��@?KL�kǸ3hlrÍe7���ԽM��N��ZY�f��(��l�x�5����.���y%1�G�n�H��J�����
M	��ʛ��&=������
+�+�����.ȓWEjtO��!;jo�i�VO�osC��ʺ�M�\w�?�^6�`Jw�q��J���!z�K>��w6C�XS�HG���ٰ��)�A�XJ�3g�`�������1)w��˒G���ʔ�6��Ė�G�]Q�k"�7,-��o!� p�v��Y�:z�Ae��𩈪��1�/��<��5>Pp�o����!��Υ$A	�L�)j�E[M�1�_\�덌��<�����=eZ�����qB�~^�;O�g���Uwp!J�o��&�k-�#.����r;���ɈtcK��lG�8Xq���5M�YK-���q��̙G�p<A�	��0�{ ��uEZ�/bŗ����*Mͤ22;�w	����k�S K�o�[� M#��� �B�W`f$�z�Q^݅�;95T|��:ŘX��i fZV�n���Ag<���PAiA�]=&��Ɵ�6M�n����Iz��7
RR���O5�ׇ[��$s1����k|����X��_s>FQl�{V9�o$��R�sW#�-Ʋec=��2:�1NT����RD���Ԙ��ٙ\UT1���&P5kX��b+W9��b/�-X9���!}�~}&�
���zMi�8���`����Ф��X\LS��eѸ~���n:�>eT�@� OQZ�
���@0s�?���[�A�괗QS���&~�nD��/��L>[�(��
��1�M|�6FVyA���ݔ��w��X�IO����Ӕ�l�Ϛ}��!����Z	�]�{3,�D �E�c;cn"��&�j���sa���`���?k�q�������@�y�Eg���F����Ќ�Ys��r��efm�h�̭t���<7�6������۔dQ�?:�]VP�W���B�i?������(�>-�p�p=#$�.��ry����j[W�Ī@�C���;>��t��/�(YNz�x���#����Q慄ւ�����\��	�֜��|ǣ�H
B��ɶ���8�O�6b�x�v�f�8���ŧ(3����T�1t��ߠ�fx�Jh�Z���%zc��m6Ӯ�R�C�c�tB��Jz|����������ٝ*7;>��S�īQ^t�Z���oN���,uΗ(ޮ�-�W,��6/<
]����?8��1h�j�L���O׀����,��}@��d�to�5����3=�0���}��i���DUbI�<>b�݇%?��O�"@_����X�;���I/Sݠ�}]y��h�d�x	�ͅ5m;5�����yϱ`�1YV���������|}e�#ۺ��_�D�3�+�mI��zh��˝A�5��Y��o� ��l����7�K�j�������J�.s�5�pQo�DeR��Bc���%����ޟ�����$��U�EM������� w �|'��ʀ�����)Z��N�h�jdi�c��]��χ xZO������:�]��U��J�=5anΐA�ͩ�aB�j���r�s��G)&��D*��2P�C�B��w`�
�Ӯ�2Vk���̆�D}�|��=��Fׯ?��Ա���`8�L���������fs(����33rM2<z)L(S�o���׽���+�w�D�7�<�����CZ�s7Q���)�+%|{��v����mS��,{����O�U��̗���,�z:_H�ꡉty�C��I��OQI)Kh!�:�PU�ʾ hS��֛�n~��%��q���U>D��^����z:�Z ��;}Q�}a1�n��G}튇7D~H�5Xh���x�C�����9��w�v�����.�|�%cr�]�]����>�A>��fD��J�'p�2����O��(�Op���ւ������J-�|SY�zyq��ύ�:�Vx��Y�o����5����6�K����>��{5z'�`p)�L��L����r�u)���R}:��h28��&��'=NJ���ݯ%$��Ba�)�#Ӎ����r!풪%�����K�*������ o+�U�q�0``dw��r�T�lھ�%c��<�]�R9���t��� �G]�R��V�6�+�X�j�nՑ׍����]�њ1�.��͞�p�~oN��y;��>��>�l�GLw�����	'.�ӓF������E|.�kQY�5����d��	�M�ھ�t�c�j��Qi��C�p���J��wO}Ԗ�_j��}��)�_�X͞^MШ����\����./�V�;k{�¾h�g��HDȫ0A��]t��U�2sl"!2䘪�1���
��:N����8|��j.k���'����s�Vw#5?9��u�t|����D'�C�⑺u�h�A(�%�c ;8��1]dTm��hp��e����^���5����9�H�7�wSf�$����@QZZ_���
^v���VO���j�n�7X\r�I�3�݊�sz#���]��P���gc�"���\���n��8�g���?���Eo����J���zv2�:�$��8P�Qyo%������D�Yr��h�-�i�Im�N_��SG��)���'�:���Rhhr�ذ(( �[����	��d��&�7�8���cߩ9�����QH�Q\=��K���d��$pza����s6>����/K���	.���[G �#�c�I�h�%����$��b�3y�+�+�G���Ԃ��$a�r���?^NkeY98ۨ�ŏ�]v�lNLK�d�A��?\�PM�6��ww���Ip'��ݝ�Np����5���K�{���W�Vm�L�>�Ǧ��`�T������(}����b���l�]�N����֜Ϋa&8t�/�I����+ᶾds�����3��[����
��;�;���N���+�̈�R�F��+�jx!�x�o< ĕ�H.Pp� -a��q�>��ۖ`�[�n-ը�,�_�w������;�9sa}�YN���hYٴo�̙9cN����y�/����R 
�ΝT�h����%�m�5T��Ei/��^��<��U�����b������&��~�7�g*X��L�P>��K�I��h��"��z}���_of;<��oC�X�Ar4�9���`jr2�|?��t�P�����|Ůx�mߊhÑ _NF�����\�����z����z'YA2ޥ�u��G1͹�T��R$P���M2u�V��	:}(oc,�R٣�]��a�x�T�B�q�n
9͈@�g�$�ݢu��]��=�����ݚ����T�'WU?���� �ې���.�6���>i�s���4bɚ�z�7��v�U�T" � 3�k(G�Ӿ��&�kn#���Y
��P����h;�w��G�t��� �E�탚)S����?G<���}���e�|�U❗t�	bҎkG�&�U
��<d���`�V<Jb@�%x�k�J�ɼ����A^���;)NH��7ӹl�k��ز.<}
����{� ���Vt�t�ק��󉇟
����_
w7ԾU5ѝvy���H��Ǘ����p腼��N���3� �
�h�X/��tw�4ެڿ��dG4�$k7?��~^t8!�[�L��a�k��"F�����B*0R�,��)Ȑ��Q�u�a��袲PY�R��t�@V 1S��'�(�vZr�L�N��-�o�g�,"�	�e�j��B�ۊ��Sۂ~0@͜�`8�M���>�Ha��E�eTßCg��K�[SA ���'�h�|Z�>8�omwۚL7i&�o��li��mn�z�>L&v(1�ʚ@:�R%�)c����l3��X��rũ���Gk�P���>>�YĦ_��T�@_�F.j9`����^�r@%�Q`��.��ѵ!���+M��\n�c���c&�ˠ^�R�/�$�C�� ��`\�ޣ�{���'��{}�ϐ������\{6�@-���8��|����>�*��������F�5���Ve�h(6ٹ�ĐY�&�@L���8���⨆~�\���.���aC��n�W�B��|26���l�ޞD�����%|>#������ rK�@cGs�x]iN�T6���FA��ɭ��O������E�������dn�ZsjMxV0���]�,Ґ�&����NU_&7a�ݢ��!�&����/�?^.�l�.8}\v���ˠ���ͥ� m��9,�5�Y;�CƦL��|T�#�(�����a��ڈ9<��{�4��eR;�~�);ZT3�ׯb���� �G
�u�3�Ɔ=�u� �r���]�k:�S�y�`�Z2Z�f~�_ێ�h�W���z��,O�Ý��Ew���̳������h�ڿ&�(�eO��gk-*Y!1��ٖ�R*҇F򰴔N
��_'�Y~����K]PR�_�#k�u*K��
yS�?_�f� �2H�x��{9�,"�6��gn����za��Br�)
���M���)�boD�uT�$�T4i�W1DBdt��~if62Ipj�MqB�x	�ټT�\&q�U��4�u�$��..�싮sH���?�AĜ_~I��{�q����V��Y��:r��v3�N�ufÿƒ_?��83Ctns6��=���}��S#�^��,#)fMb6T2��g�euI��Vev1�B�9�Ɵ����%`&ʎ\�Z��-.��,�M�~|���2M%T�1#����3d���g���dc����������Qq�ֹ��pi&!�:�M�r7��1A虌 Ƶ�Ý�����,l�j-���	�P����ǜ��:�Z��͓�<`�"w7�4�_;4n\T��q�yJi�	a(�n�3u�Xn?o��~�M�۝�\!\��jԿWm����}1�Yyk�ܭF�y�E�����Y��r��˟�b�&��(�84�����ZC�ǚ���bӟ�\�`����:���I���M��(_���V/��l2KTT�W�5�@$�(�h�OY���Q�*��J_�C�����MI$`�NDQ�NF�(si�߁Ȱ��,�/�Z���(*2����h��P��°�
��*ۇ�5���C^������@��A����:��q� �!�N��XK�ۅ��	��c�M9 �i!���M=F�mР�a��������Ba�@	��}��p�<��Ŷ���Q
�e�/��� 5ġIa[�cM�\N��
�t �������(?(��Q�/�+��O���0i�'&n�`�bV�]� 6oG�g�oH���l� g���3BE�jq#ږ�����u1�+�1'�p�`���7/��dP:��t�tX?�Qw8�W>�7���K cW���2	�� �Yy�)�q<z�.^�aL�$�G��ԙ�W0R���!@��W�<64���4���(^�Tg�x8�W#���S� d���W"я :M�� �2͹�%��ۄ<tX�x�v�z6�5�� n��$��7�Ǻh57�`h�����v�j�A����q�q3��nY,� ��rc7�jU=A��-:�36y��9�j�Yxy�"q7��0��0��98�����DN���\n�׋��y^T��⁐��)�@�٣�h�����������'�Z�Mqi����P~�N���n��}�9�����@�b�|���rQ��/�fs�qa�ys��L�3F��P�b�[�%{��N�}����z�XY��;��E���{��q���&(��O��MV`FD�޶�{o�2l��xN����x�O�6<�uU��{�����e˟��Ou>'p��}�`9Jiy>=���Z����"!߸����#��D�⿝����m����h1>%�a�ޟ��6�$C;�ھ�� 7P
'8v0m</J�^�W�#'��K�å�X:��o-��Am�5 q1f@�����V���A���Ⅽf� W��'���53V�pX�j[�ǚ�y�H;��(� �!Iwk��4
��ԙ�`bB��}a�����6���]���κ��KM硜�%T��d��u
*k��`ط����Bt�Cy^GlYY�;ᯏ�/oG.O�g�G��N�2��@�'���CG��zn��u͏.ô�]R)�˦�����eca]Q�]�X?��Q��;oJ�.6� Tcr��V�/��t��YU	�Xe��jq��O�ᯞ��yY�0ga����������
�h7QA�Y�-%���!��.7�#�[�\���8�8^P��c۠T�8Ý��d*�T�����ݖ!��\��b�H��}�1^^��U?݆�ubr��`Z_����c��-�m�O�!
�Еￕ*cA�f��QKs'f�[y-�R��> ��Ç	2�U�5�c��~���b��|�)�G�L�����h���-X!�ƒ2n�0{��?$�s���z?'��i�XX]狂��6��e�]�:�.^7�f?lB�p6Z��6(��O�y�)�Ο��f�����p�Ѿ���{��A��Vd�VIvB�%/9i��;鮽t�p�GQ�L���/�)SR5[�������]��Q��S`���S&��뀫����b�5�%�"bMض�Q܁���E���ع��Q���id�!mr�ag}D���X���k��x���?�d�}%�>��"T7�r�A���N���χ�SUG�X~�q�T;�y8xrySD0u��ZG��6}]�=��P�ӳ�+�����;�Dux+	���l_��!
�3������.?W5=+�\�t�6q[��N�9���?�0���v���v?���j��h���j���j�߈�`�W�.stf�/y|�Aq*R�/�'G���9<v��Y��Fi�6�;��&"5;=Н=���_��wژ�	nV�`�'#�O'�VY��߮ZUA�ŌQy|�hu���Z�h�o2����j�N��4�� @��o���&e���'�����}x��b��ꞓ�LPw*^����L�):i���M����;]*�u�$��*3z�7.M�O�ȹS U8Y )2����)O��x�f�E�2+���k��ꔄ^]��ݡE���K�U�&��=� ~J���u���5c���^���ӂJ���6�	����I/<�;+]G�6�Wmq�ko �_s��/��E9���<6NZR'��@ax��ǟEK5Ê�y���dO.������~X�IZď�n��Q����r��;�v�M�{8��͜Ų��1/�K�p����$�痀UY�S��_XL�Ȓ49�zY0����6���F�P$����2��ƛ�QN��Y$/���^l'L�l����^Z�N���	�~
��|#���r!<[ja}|�NV.�ˊ�H��SD���MT�:e�0�O��4&W���]j�^zf>���c�˘������6�( �i�mp#3(��&�O����̈��l)�P����DK�b���
鱃��=��ND�tc>T$��j&{�f4��jB׶�!Kp�����>�Z��v�4sʛ�Zz~ځ:�Y�Q�}��`�|��%�0�9�5���ȷ�d�{Tp�괕j����d�P�.^5]z0#6a�;(xBw�#ͷ&\u"��ڡe�Y��Hg������44�	Z���*I�/�x��%N��傢�w�'����i��	�;�AT^s~�����h�F�Kp��ٸv������GX�%;i�
�ڵ��\ �����]�VP����+��e���l��ͺ�ł�b� �g�
�	m*h����e��sTG&r��-�F�Bĺ%�|5��w��P[�HEJ����ƻzwHU����K�x;�g!�Ì*��ݑ��N���|��h�׬�jB�ྃ���i��3�{q'���o6}��r�,��Q��[jj��*��M�%ԁ�E����� ���C�Ksر5��9Fӻ��He��ޓ��hu�k��bo�͛���|�щ7�.JK�d��N����8����f�H�.�f�B�[/����,Ka(�Bz¯�m5���8ۿY�n�"��&�j]3�k&�b���J�J�W�<Y�%eyI'�3o�$��e�L\�iD1$�}�y����tC>e����k�%:��؇ƴ���_�����ݘ��X>Ƴ��&����r����(��]�^��p����X*�y�.�Ω�q��W�����xE�����W�T"��?��BxT/����d^�x�b�% A	�����`�LA���ب��d��N�DE�\����`��0S�Qf�ƍ�cX��(|���G����U+s��u˾�\F���y7���3WE�]���0�d�gu�M.��J���F�}�J�>��(Y��?=�<��W�����j�ޅ��#�0l~�떜^uPTn��V�
�^��y����]D��o/1���;��Y|���/���I��(q��^��ZGp!/h=��ͬj+�~Z�B�TO�|y�c)Ops��p�%�:�M����%��;��ͫ�L�֔5d�L�������|,|�꩷Fc�!H��/\ډ�7C�̈ǜ��Y���ﱅr��'�ԯ��q�ycl-��?�~2��<���3P��;�whUµYĴ�]E����B�١mM�g+���Wu"�u)l��=Lee�yX9z��##sEY�Lӟ�-���~��54z�c0� z������Ji�����fi������jn��?��$PPz�6t�ĻUO��/����^����׮bMz���ܭ�N���U�fF���i,�.�$�Z��
<�F?�����o��-���}O��퀘嵭�����k�]���6��w��؉��+|^�QCe'M�S�>e2#vі;o��}'c�n�]5�����;1C���^����`�l	T����4mm�؆.mK{
��������I���� �}GHy��r���|9A���N�[
ݳ��8����K��2�e�ڄ�<P�.*�xb�W����Vr���S����]�|k>�r)��Ţ�r�x��.<?̍?��'�x�jƌ��e ����~��I��"�o�H�8.'���۶�����u���c�t�pү�ɐ*��S���;��l�}���lF�+���l�]A��۔�\����۩�_��QVD�������t�Xלs<�/��<�,����Y�~��>xT�����Q��_Oxm/M�����Z����&$����FF�0+�[Nz�7	T�Xv��(X��O�,�3��,=/i����T��xM򺡵XߙTd~-Y~��	��}����uR�
��p�����kl�9�U6�̌x^���-��{>X�Z��Wq4ѸЧ��u�jс���;�E������x��Mh��__
Kz'�,c��wrZ"�`�6�Ƴ7peZ�o�tdeȄ/hkJa�KT~�6�o���7�������ڻ����`�ɿ���J�9������ۅ��۔e1����9-���1���y}�1y-�5����e��e��4���I�C�@��yo�"��G�"��i��O����ҥ\4�ٿָpXN`>�@B/hH3D�.���}r;�5��	��aK��X�Y+ ��*���i1�ݗz�qĮz�8���Tp���n�,��'*�O(T�K\u�
D��%�H4�njuu�֔mU�,r�g۟��Y,��hO�;�B6M_^b�t�g!��;�P��-�z���$�.,>������x*�jzpsD2��T�C���Y:�y��@kUȒ���:��k˹���zd)��ok��t�yW
,.�v���|���ꌐ�����+m[À��*��I����"	�������ލ9�/.;�9R��JӔ�Y㣨�a`+MuyS?|2B�i�9|�K_���XLZe��F����~e�2X)�1mª�b��;����Vg�	]�S8	r�/St��,H��T�e"��-�56W�
��7/��o��[�$�U�(F}\�bL�B���
<B��K!��g���,���-i\� ��!�Jcq�T �w�Ŀ�?�!��\���CCi�Z�,�r�)S�<�����in��P�zw��|�}͈),O6����,�~y0��H������^*���� g
gƑO{2P-����<nЌ�ա������5 Uk���3;GFY$�����7�%!M�h�5�ܗ�5��{LT�*&��Lw�7�&pj�}�ͳ��?�x8�)����-�L����ū���8�j��a�=C�xT+���~� i83J1����)�ҳK� @|��M��I@	�fA��r����S5gHN��z����D��)���0�z
��Q�q*(�D?���~�lV�O��7O�=��K�v[�$����L~�Y�1@D35@}��'��7���? )j����fp��kh��a�Bu��`�<��Iv�����
^>����Kވ򌦗R��1Y�G�T����H�[��Q��~ڵ�d�"�Mh�S�>��cŦ�eE��S7�D��F��+��,�������bie*��?�-�;vw|3�@vO������_�=윲��@��,.=�q�oh���9%I��W�p��w�`�2?��,���^u��.�Bʕ?���n]S�����(�7�G%I��c(�[�Q1�Z��u{{�G�Ν�`[m)(��A̿�&'0��D�����A�+g3O (L����t�V{=����S�d�-,L�h�f���V^�0��V$8�=g�Bt�M�e����?���޳R������>�J�mF����q�Z��n��Q�P6
�<+�{d@ÑF������%�H[�PeW9�'#���]�%�3��c~��&-�S��6�s�A�}9;'�����kr���U����
�0��n71R&��U�TN8����A�ԁ��Y�e<�'��`*�SF��FC.�:e��<��<nd����D����yB��1U�d:�J	�BZ[]>M G��`�z��r�����K�������ҦoW�Ar�m�烱>7p�[��X}����R1��0D~kU
c�C��Y+�����l_M$�Yw4:֙�5��)�Z���A��21c(�`�V�I�5�K^�%�6|��P(S�q�}�-�h6UУ%/G��b6�o���B�z�WA�����&����x�|]�\:��C��Y���ڣ�v�R�B�}k �����:B9Q�C#�v�LnP97K
���ڐ'���	��H� �XL�i�ao��!��}z�,�GK�=��:��3�� �['T��I��
����i�ې���1���PDq'w�@t��1���	����O����Q_�
��%<8��1q͌a�g[�#ƀ�X��ԧ����tE.XCW2��/w2���d_�"E���|�EeNg� �D�ŽD\���]t�!�������]J��Э�j9��u�CK�]��|����
6J��}�m�$-��m�yM%uBT(��6Mtn{܃�XZw�7?���i��)�֎/wBx�p޺�0H-4I��b2�kOI��/�N*\��?���Ew�NB $�`�-Q-�����f��c'j��O�r�+�U�3sj��zT#�5٪�P��Ũ�Å��S��v���*_܎����AN�P3�����l�%ku�]=_;��$�
���z �A�Cn45�� �ǃ�|#*�����J@Ir�O�"��Z�Ѳ���dKC�I某�%�p/|�žJc�L|?u!�� 7�j�	B{Wx>S&g�ɟ��1��#{w�2�c2�-���(�Yy�_X��s����t�jL����0$(�0���5?^4x�M��J��j�})}=cH���kCdK$�-w"�	r�ñv�]j[Bb/�z��Vg̲���8�L�ispk�¦n�L�8)�����h���J ʅ�4��")H�eHX��l��m����L�e������Ӻ�s0��������7�\�B7��
F�C*hރ�����PCg�����]3(����ǉ��8��r2�ڕ�B��bV���6DT�/�=�+�V&NV��@���w��.� �C�Nn��Pִ�b���=L�sZv&����@����C���݉E��d�g?*����"z�K��xg�Î�%��T݅��Ϣ�~ ܎1�/��s�4��ٺ#n��\�G��W.���߱�"��e&'@�Y�Gf'F+�����0������(�gr9�T�Gm�;�{�fG.c�\�N�"j�nn�%!f�������2T3�!0�8��=���Ϛ#tbq58О9c,"5QqbA�S_4'D�M�{!���>�#�8Z�rWn6�<3�]��{��Gf�;|�b���'Fڷ��CB�%���Ɇ�5ﵵ�y��υ�De!n�J#�~��%P�D5��o�� ����g�,f��Qq�Z�t�_��d*���EX8��KhN���K=
\Ծ/s#��#ip^?�������B�G ��(���:xܕ`�:`:v�.��A.��_+S\�a)<�Q��Ԅ��\CG/�}�ق��9�Wf�)"L��� ܲ�X��/��*%TޝZq�߱
@�dq�?ŗm���#��@<�Z��k�kw�g�I(��4>[mݱ����%anY�r}V�V٧���K��@���U�����C��]
D3E��7��T���V���2GBԎ��[86�A�V���..�n�������x�S {-�DG,2��VM�| Mu&����*ȑ��H}�u�n���=&ꐂD�@��ba�K�M"�?a�S���P����0�v�)�w�l)	��a��)�0���u�����K����9�ޮ?|:��U}�x8��}N)���_����D��$��c�|�vzp/��j>��o�[*7R�*�5rT0ᴝ�.�?믔���3V�*����%8VUJ����f���9"�oz�s3m�j���� �{�����������	nI,G���98��fG ,��;�AgMP�=��U��<R'���!�Aȫ�SZv̩�ԔI���1`�l�~h-@s|��R�N�j �C
S�tW ��h�oD��D�=�m�����xz�gơF�"}�G�z��A�|6���R��ۺ�O �wEۘ��_�����i�n PL�&���R�^�=��?�*j~@"	0�UV�WB�6ħ}+����)�b_8�6�� \r���>��v����,y��%'n�W��z(kh@(��ť]�{�'��g��I��j<A		}����`�u�S��Mn3����s��&�E05MӰS#�F#�YLxdi�i�s�#�w�|z�0�&7�NPA�5Žߤ�����qy��k��}������2UtV�J���֣V�d�U6������˔������.���2�Ƕ#7�c��EO!ӛnlkty��k@`]�q�d2fF��(}����ʡWxu��O���EjyӃ�|
���R�P�%o'�Eܝ���}��{v��1a���}��P���(�W�Կ�۪�Ѝ�ܖsmM�q����$��V}�Z����c���Ыv��P���\(q�L�W��U;/Kq}�����vb��#���3ި�Y$A����+�U�򜣆�����P��7j+���Z`*?G]�;�V�!%�{p�ޭc�]AA1*�ڍ�op�՛��+����!7xD�<�w1޵�p��K��z�����.0
=�7&{H��n��IS��s���=/g۽r��8���������.vC�и#�	���+[�=��jqC��(�#3:�aB�B�����Vj&����6��^&QM�T�ϥ"b����Yg1T5T�Ŕ8XO�EP��m��b��r�)O	6��X!����A\Y�6�f�(��k�Y�a�oY��"�M�X~�Z!���}�w�	n�V'��� �r\��Z7����vzƴ)!��6��aN�L�N��zI~�����z��ٯ�ub���fDaBX��;C�@���-�f�^sbw�ۇS[,�ޚ!-%��5O$����,j�y��#Pn����#��0�K�$�Go]n�]gi�}o �*4�ܟ�I���S���c�88�]�4���L��	��?�|)B�q��*5Ǝ���b �JUR`���]]�7��[_Β��!�)��4��������w�s���*8���m�b9����������K��W��kl�ڞ��=�ia�X����tfkjB������u�����y2L��cߣ�uZ��'i�e҃�r���f�~K��a}��5(��H�����w�3���!�H#2?L�&T��rw�p�Q��LBB8PKݤ�L#��
�Bf}�Y���˷��A|1�4�mw��w�:ѷD�g��͑�.7�������Kn/Ab���a��)5J\P%8e��c�d닯@�.�2 �]���8g4n=N(J��\�]s$\|I�<��B����\J���"G0�ln։v18���s&�^��������ڄ� Ot9w"9n��苽���c�Oޚ���Cu� c�v�B8&B�0!ב9��~��^��_�q�Z9�ü�6HY�2Z�Z8��:,'м�q4�d������)z�"���W^��C��(������o_[��E3�uiב�k���A>B���v�R����i��Җ�װ}�6~���u�����:�OG8cwtQ��\�T={ʬ���>���D?����3Ӳ�:A/+�q���֭j�\���a�t�n�z
�L��Fi��O����kԃ����������AL�E������nO�ܑ=��ҕ���u݆`����,��yǝh�G���:P$H�T�,��hr	��>P1�j���тe(���F�x)��x-�N�{��~R� @K$�sR0�MJ�8�ǆ�@7e��c�"��LØ� �.�k����@��Y9�&%@����w����:��S������]Xkt�Xl��:"�<�<�z���}�vdd:��nl�Om��2�v�E����<����eGh�u)Ռ�����n����R�w-�w�%��RJ�䲥\�|���x�W_u���o�;W�4��� ˃� (���	��ghG��@�]P�����z�2�8=��xyW�?�R<95�[�+ڋ����_��s���q�}z4q� X	��5TP���������	�q���F��1����K�+	A�q������͛�0S��1C@���5^9�T#��ۇ$���!���3���s���8tn:�v�k����˴r"��ͧ���ϊy%;��,���ozB��D1n:K�L���N����b�q����-Y�EP�#��1w�=O��Of�u+)���n����ǎ8�=����_S��r����,�Ӳ.��:Oڝ�m���F�I,c�@�|�$4%I�����`U1���׻t��|�ھ+�̥=�@&<2��v�/:���| ����^�3����; ]ͪ��<�b����3���^�����xL�`d�r��c:�9Wg9ƥ��FQ��M�	NB��~+�����ig�;�-Sj&��^�x�}n2(���=;�(�v�%^o��X�$����S��=��7��@.ݜ��RL���m�jG+z ��i�Х�$\�B7����s�@���5�׌��|3��G����,���>R�^����ł�A�*gh;�S�iP>�KCy\3��q�Y �2��T�@��}�a_�!ۛ�t/��<�ܝ�:滄s
iLn5��-5��FP�v#�HN�I� �����Vxw��i�`��²<�'�+��m�EÚB�<9b�ऑ�c����`yW��"/���$�β�Z<v��.�mVX��A%!REk�n@2�Ab"A�#�<��2^�^[��d ���O������ڸQĶ�UΛ��	���p�ݼv��������0����B+���F9Ll�8L�6����#32��oU_A�
�w�1�m�04$��;�篞v�GP �'V|3rp�����^�*��16�_�!����5�%�t���+~",���pQ�g3�ytE�E�"'�\�Ѹ#�A��qю6dJ��K؜Y�-LTgꧣ��)j�Q�/㱣f��}�
�_�o�z��ۘG
�u�dĹ�β���bێ��wo�Ce+�O#�������>�͍�Y+Z@�nB��$yL�-�FM��|��D>@�F�O���bW�ڔ�g��)�.[�ZF�.��7nù
��|%�p��9�vz�>���V7ӵ$��t�������ɀ���ψ���2y7MY�!�((����'�曅 �����t�����y���eE� 9����*>�R�M.�-�B#Kа��i��d�y*�Đj�b$���
���|3aF��G�l8��@�{j��z&X*� ��[9��P��
��~/�/��<�� HL���W�9X����<P�P�������.q��G@�I�jr\���|���n��j��?��1�V'}�C
�C@�1=��06��
����W�v*e�;҂з��-pr�i�;�o5��ey}���-�>@T�k�p����
����V?�ّ����124A��ڣ7y�ە	��c` T	3&��!��G�#��p<���P�������M}Iq $���f�*�6C$-����O��`�OܜI�vyk��tc��+��ܸ�X�v�����+�ҒR}A���1,�8'����T��?(�~Z_K�j�����X	p;
k �>�ǕږlL��0�j;���Q[8����G�2������ S��NAVR�<�����
����y�7n�5c��+W4<��b�ٌ�=mK� ��0�ҴЂ��BR���_�T��>б�a�X��Qg�괔���Db�K�@<3l���6T����YQ�2	��g��ĥ��K
���v:�g:~����j�l5�>C5�ﳬ�����oij��Rl�l�i�p�y��L����^���}�L���d�Ӏ<7~��b�<Y���t�xT
��uC-�Y:y�QT�<�X�`��7/�L��d�?�GXL�|f	p���P��m���z�7�VfҸ�b�=���c���`_��xr��H�po�+l���i���ޚ���XH=�C�_t��D�cP����.�BMM�J�����aO���,3�+
��7YW�F0L4gn��;��
c
n-0*��xTC3	f���I�x �=m��\�|�� l&J���/v������֗������>�a��/���2��A���jВ��
~ �F�8��h~�C>8mu�a���t�Y~Q�q8nPq��A���	�G���A�hŊ91��;�����~(���:F[���^ۯ�A(*~��CЁ`3��3-����u�Et��kA���I:�C�wE@��m�vaiv��:gv<	�vFu���8k;�ݹF�u��c���GV�iJ��v��a�e��?��aM���0��ޛ���iV����
�zh�U���SUQ�5���b8�P���Ga�l��@菕��=�a�T]=��r���3awww��f�g���;�Ƣ����:������b�>3����g,n�hʆ<nԇ;ԉ�;����q���/	2�̰P9^���5�Y��A<� ���wA�,���6����/�74>O39�5��0$^|ߨ�y)>o���E���f�'��ۨ�bZ�h��C���{r��P�� ���b�yl��{�^�� >��7�ׅ�����f��qes�G%p��mGp �6v�TYY��M�������dw��|J�!')��|�zP[�����d��/)y�诣���DE�_F��R6~:����`���CU�m�Ŀx��.O�'��B���>J�]�]<�ĖO��J�	��f�kJ�E;�i�� 	�W��B/��D_�x�.Z�km7��۵��rVI���\U`�(�O���|�[��/6EV=�+��v��%���ܢ8`L�+�#BR�1zZ �"T�I~q��8!�5V��pi��38q��T�Z��Dr)���Q���s���܃�+m^\yt-×�lT�ч�3�|ot8ZR5�bn	2�%`��04�d�aB^4��{���U�T�Y�,�E�S�P?�/G�&��iq���j��	C$H�!*��s?P2Wr2vr�n3��C��SX���A�ik��F0�R�� ���)����G�Oh͑b�&��k��ς��E���Hg��H8
O��Y��a@��� ��j���C` �B��TJ�%��I���$�q�Oh�K
���?!��Nh�?�B�����{��܅d��Z��-
+#q �y�s�Phm���a)�`?��y�?��OB�lSޏ���s�&*}�5t�w��"��?�AS$�!���|�i������[D�jw����?6���UW�̟���k�L�`�����CR�[42h�h���Cⶅ?�R��2�5$��!3����ꚊH��G��(&�&��j�'f�)#K�-�&!���B��p�8P�~l�����~� u�"r��\�ȝ���z�B��7��JU	���5'�v�[ag��ߠ����
Q� �A�4�R�!'i�Qg�p�� Ɏԇz�N`i��Y�d�Kի�Iq'�P���M��Wq5�EC�P ����H�
�C/Ifx9�ǒ,V?@���=�?J-�\�>ް"�b�'� ���5�(���c=)zڪߢs�A�̜t�(XQ�4H�Ұ�����2��-� �=DtRf60K������#�}H
�M]i�/��|���߫�������n]iW�}�	_��t���,l��b�= c�+/L��0�!,K�� �� �H*��hPj����J_���s����M:�&ް�[0��A�x ů��6V�ǩ�7���Ö;�o/ w��/2��#�#��)����%W:��$5I1��(j�!���Q�@��$�u=��?���j����u����\l �o���l�+�
������T1�� ���ΰ���Z��[���_]�v���o�3��z���(*�@�L]%a7vR��*�;���7K;��}�ӹ��~)�R�c��[�W�WB�4[f�'��*QE�q�[�(wȮ���#�ז=�������v�7��TV�����:@�����(df��ޔ��Y{���๸~��p�z�y��+�avG�4�U���!��-����j�]��dg�>�B�Sbu�=>ڠ�>\��j1PY}���2u��;#u�쑞��<�:�x���q�:���l�Wj%R�{x[�^�ȃ�A�n�Dl�|��<��%O��\��u���6I���8$!��L�J�щ����u�_����o�}#<}}& )G�òT�H�q����ڞ��|2R�]�3�!��|����g����(Dc���!�	��q�ߗ�h���N�t�/�'�����EB�� �I�����&�T�5�(f���P��"�B4Ht��P�:25��ȅj�#�M�~�^��ܱ(��NC*��N-S5�&����;�m�������f��[w.�~~p�(�����ŏ�����3��A�;l�x�{Ux�zg�\ʱ�%�g ���}�O6��B���M_�?Q�������[t0
����PT4a�hڔ���������oF�2rrv�ԛ�㯅^�q���Ǔ�����j��ڼ	��t�HE�ނҫ�J��(@jD�H(]@�H��.U�-�*z��]��7�f��53��䞳���쳟��uW��E<��J%�И����rC%6dA��{�f��1�E�5m���_ד��Y�7�����)��B]g�O�b/��)���yy�&�4bƋ~U�Hs��uE��inl(���L�jt��`��N��ht��n�P����W���a�雥w�~�JV:���m;%�mB"���R ��{=߾�,���r����7����c�V�,kC�rw(*�e���#���v�F֜�
���^	��g�?:bu��;&Ism�U�f�Tf�fZ|�]ay X�3����>���޹���Ns<�H�d�@�m�s��Ϻ>���|�~���i�5%�s�hc�k?T�v���eH�N\�0ְ�[�im������6L�!�$,Z��ɋ�f�V06}��S	��3�,�q',���:��jģ��#���J��?j>3��_B��t��*�h1{�yI	���T�ߏ��2�kJ�"�\O������_�81r�k>=X}�C�)��>J\g�	H-2L��#�`�V�IǟCIqd����!��6����x�X1�8�*���1�dE� ���^���X�J�"��p-�N^��*��%l�_��ʇeo�^�to2<�����uRVs����\�[qO���m�̗��>>2ҿ���P�g>�&�(�_���d�/�Y��0ik	g���)�
<<c���A᎟-��L�����_{��tv�����;�/R%{��^��ף>�U��W�,���"�3d�{�²�?,9�5�Ɏ��
�O��̴�&j�[/�J~���ݏd�-2"�ʌL��#���X\��~�M�W�-r�#࣏Qq���VT"զ���d���h�R9@R���ё��ExDu�u�?�ѠN��9f-''��>�6��Bt z��ӫ�(�
��틮Y�AKE���.���鞲֡��@k�U?V�Zd1�2�$wW�-d�@&�A�\���A���hSI'T��C�x����&�NN������IE4V��J��JD�Pxj�7�8�^[�t���%:��!Q;NO����;��@��X�FQ {�-�w]p8ִ"�f��[mS�jW�l��Y��#��4O�����j��
��g^T�s�Ʋr�u0��7�\�Օs?|��u��������f5�Qt�E���OP^O+TY�k{~4�|
�#㝬��M����p~��HT�e�_��V4����'��g\N���J�|��do���*pNnnL'038GR㆖�s��o������������+/(Rh��z��Z67_21���6��5X�̙�݁�#�y�@D���P1���@���� ���%��a�D	Gwd�EX�)�1�/SMw;�>��Ԋ���=LS��[��P+ d�95� ����Ŭ��z�k�U9'�0KY�hW �Z).Z_��?�h-�D
�BRr��L���q���n:G˦*"���
XSu���%�����nB����o������_�#Da>�A����(h��e��J\,��E��"�ח�>0+��o �#�[�q��B9�Z������ 0䥮W�*�!����;Z��@�:�O�@P�m��y�0� l�#�/�0U�DH�Y�E�_t.#?T{Z�V�L֗��9�1*��;i�0�m�����'�̽�<v�T�ޢ���/4Є�Z���J��Vkf9����FI�T�ԙ]Q�0B��N���{!�6q�vƻ�
��O��C�R8�����Z�	�Hۗ�u|����"BZ頚r��i�v����ɩ�&���`��:c���mK�0 �},��ϖ�8m�|����a�ʳ�'q��$�W�RG2��&���;�|}��� ����r6��J �X�2$�����R<���!V�a��PI���{M�Fu�٫�04��+�\��7� �_Ri����*u����'�Y�,���"�Yp��p~��6vvvi))���S6�2>Lm�w�2���)����2�2R����<S'H�T�d�
lsC5�4��?<�6���`?+�4�(X_�[�l�k�iZq�Jz�V;!z&�+�����m-�2Rl=a����𺵦'S��9R��btuQ�t��9�/u|"lgR'�Z���_�±�+V�8�D�h%\W��乚&�7�mJ$���;#y��O�z^x_ 8��y{���ADa������.��x=���D_��*+T���07�5e:��>N��(�][�˾8��ୗ;D��0�����Y�8����[�˞9�����q��G���b�ǡ��2t6�<т��`����x���v�>R)�k����'���/����#d={��m�Y	~�b#t�h,��.NK�V�+y�YC��.w�NYT�kI��>��E�)�-�gJ�.Q��B:BHG7��n�s�����/^�s�].��;�@�Ҳ��g����Lwr�H}	�1�� 9fC
}@5�}��i^C�^�V���q�#�9�U��a��~�O?�
jw���\��&%��z�	�`�$' u��:�k.^�׹��{��>�_wڦ#*���_��g-Q~Q�2��E������z�m������"�$�S�|�E?�h\���1�z*���.�c]?\]s:k�J�/,P���S3�_�����_�ƪrEB��K��}&sR� )i�Fx-q��N=D����!AEت�il5�Fh�=�[͜/`�k®�xX
���7�0c>-�{��L���[��m;s�S���RHŠYg{�۷��0�������t?�6�n ���X5U����&���n<��u�r�JH3ou�˭wM��r��%<=+7�C�ۮ�Q����rj��T�|��Y)�N���*z���Wz��Ol�}�~6��W�L�2�{����j���(�d�HY0N� ����C�ng"�Ķ��iХ����j*��ZFfl�	�C_��n��A�6�"$5��!�K�1�z��)�;z%�^qj����b�w=��d�W9]��<N��.�,Y�?N�n.������O�"��3�fl�B����.�2*$���T�g̕/�v_J��?�jI,[e��{w-kǿ�p`���t��H�ÖN�p�m�g9܂-F��2��8�b�M��� �ꛗb���չW�'5ԛ�NW�P�̖y��&j����p�7��p85���[r��$8�֔~0NC���H��k쫇a|�yee�1����'F�]+"�x#��zJir��b�u�CS@06��4u�*Y+�	.��'��ƦE�VO����^]�*C�{2#cS<X�Ɔ�j����w&s���Vz��eE�R6X��F5�g�BU�t)۔}��0{�)�&p�,WEP�tɧ���MV$�΍�2u�8�������\��;�1��𫡌f�J� =�ɒ��w3���W;�M�b�*)��H��W~�V�I�5�O�{���;qx��o��P��锃"����	�A���Ch��*�w�Zݭ�^�O\��dx�i5�;ٛo�ہ�q_����Ę�N{�;���h�W.V0�x��"�v*��ʹO�5n�������Y��	/Y,��7���ke��A��ƎW�]�7��/��)f�Z�X	��ɭ��5�"�j����Ki��fY2D5�ۯTm<v��&=ӝA�m����cU���y#�c��8�O{�^w $��l{�@Hh��0�o�k>و~����2gH+[YY=m!��}n��m�7��F[6�D
�Gp�k�/�Z����ܳ��YJr���8U����rwj�b=cyw�i�����qc�˾��?Dpu2��JC��M.��ޭcA惱�ic0_����+�_���b\g6��:_SC.�,���!Q�]''��i�#��n����>i%���L�%-A4�����V^'L��<"\��saw탹��_��>/,^Y`�:��069���Zu�5;[AA��<X�#:��<s�������#c�����W^R���~uV%�O!
�j��K]$�>i�d�U?z^�����Y=�[N�RP�?ٞ���޾�>:�w�Jq�i��	�\b�����������[bbLKU`1`�v��[��z�ּ��\���N3�f�������sۛ����k��V�_(���N�a/i�~mZ��^h�x ���;�7�[��(�4���s�����M�;�g>n���舎�6��(�0���Q,>�/l�HP��!��3ȁ��� 1��}�Oӕ������L�Sp�w��چΩ��HK��r~�_��{tyZ�`�5f���Kw,�(��<C-�ߺ��.:�Ye̲C����D��$Q]^Y1��(�r���Jng��m�"�5�������ۘ�W0�Ǆ��{���_cA��G��xm��g��M{�n��o�6m��ķǊ�o�$�:e~�.6m�k�8f��g�����T��"�U�&�I7,��t��M�n��C�񍤢߷��'���ȘE(���}���jK3L�rk���A��D@���ag�<eD::J�9.]z���%W�֒�O�H�̘�1餛a;�^����5*�W�I'����JR#9�@W86��tz1�B��!��H�9:.�R�`�+���n���L��r8>"G�!��Ǐ2����F�`]�]gQ�4����ɻk�$��o۟X����{�L���./��~���ߙl
�%�������?8`D
l�I։���Yg�8�����RF��U�8�ň���{M�z�6y�vZ��b�X��;e:)I���?=��o���eⳁ��3(�Ţ�$��{��K,W��fw�d���v��@���g�B�s�㙂�tl<QT@;�~7gw�������V����;�� ���lHK���,�TΘ��f, m������,�=f��y����	�I�m����ӂ��Cb��	\?��E����_��ֿ��.{��������Pq/5.�����Z-G?EQ�	1�%�@ �0�):~�w��d�h��#f��Y��4���<fox�D������b�V�"E������&o�E���jT�b\Z������r�]32���E��-�BCp�������&�E<Id}���"Ƴ���6lT��K�z�ļ���;�4�7n\|��[�J�lp���!�AD�x��0Τ/K��歭�­:�8�+]���ɼ���J�Q 2��]��~��
�)���x�`��D�00��8���/p��^��q�ڲNu��[��{-�2��E�j��y��U�J$<+ #�VW=�q�&�Z��Y �6[�{U.Hd����%kve1���.�,z^������%�'���O��7c���H�+��·}��㶞
��ށ˖hj�ӄ#��.o֯tZR|�k�/��)#y�f��'�H@fXs��n�Ш"V��m��*�U�ٌ�~�p',����~:�\?��P���������\+p�gkP���
@�Z	��;��Ջ���@(����d::���)�R/�v��F�6m'\ھGt�q\���3�;��~�0�Dt�ot��t�ԁ���ͯ��q�r�p�M�H�g��d�~���Jf�/#/���a��ebhg;.�N��r��͠���p��޻�$.ζ��NR0\;�hbi�>��T['B���Є"�6!M�SS`��~�(����z(̋�)�Q����D,7G����`���o��JUN�GƦ��`;S�/XOqY|=gr-ѻ�N��!!*qz5�^k��9ĩ[#3(Ʉ[�8�����?b��K�<Q�$Ԟ:B�n��2�Mv�y����c%R�nL�y
�5Z��w�/菑��!/�7*y0���*�:�]������rtŚh$��ܸ�I`N
�K�n֍�t{ᒧ�e2�����K6NrzM;@�-*��ǭb`y�^�G_��[�_�7jj��1B��c���N0�V	���b/A%^9���y	�r�}`�t�w!�C&�|L�y����ߕ*Я:j�O�@0rF������(��R$�dg���x��S�A>���ڄ��y��������:Ij�ih���c���:hJ��Dm��G\���3�=�F��?b�����������Q��d7:XxCj���9N������(�H�-�%���?x�S��^���< eK��q3�%�e�(+��P>=zs�E�7Y������,�P��P�Y�*��2J�~��DaT�=Yb�m�ű��������� �(6Q«�י?�싴yް�[�˒Q��<ojoh���P���o,����!x��E��k�o1s�n���m�&ry��;s�KZ��"P׶���2UK�7,��.�~�&˫�I qs�QOV�����)�F������;���51���[�G�������6��Џ?��i�W�~/��%������~�,�6pus���fY�	:"�jl�7���7ǈͻ��G�������.���ً���<����`ff@�����!�G[!��� �t�lοi�إ��C�8e�6��g+G "�� N��W��d ��i 0 `M���i�E����n�mԄ .g���w�e�� � ��u����3 �\�Nˑ!�/{ĭ3S@3/�T�T�~������`�E0fi�ׁ�~�гF�6ZV ����|h��xuۙ��; x?S�n�O+d�%hX(�U �
=��]�A���b�
���W���+��
`y��%7�؉������"H��\���V_pOCf���JNoK�!��ED�Q��2�j��z��w�h�|��O�ue�և·�=?[�UC�R�r�=�a��+�.'

�Oߧ�A�>�������+&�����D�C�+1�\֩%�������ww�G���G>���_og���������;��D�큸����������޳����U�n?�/PK   �N�X�&�}[  y`  /   images/982accd3-ee7b-437c-8e9e-7ebd1fcbf7fd.png��W���x��,@���$$��[pw'h� xpww����]w���{��p�sf�L�tWwu�S�]���(�P@ ����2s��{����[�<�[��)Z���@tq&����醌����Q�ܕ�ã����0��Ќ�P"��b``�E��X����t��a9�檗�����EV�����*f7M�?!��ģ��JHH�`�s��m+�>=,?��8�B�ybѣo�h�I����7�.5.��}7�O�3�����1�]��fPz���	l5\B�zB���Ǡ�9�WQ���t��ԇ�t�D���=$9���y?����K=�`�?y.��d�bh�h�� ��;|4��e44Z7���A!Ɂ��Lс3N���R����BS����d�����_^��Fe�v�����t<����)^�"��y��(�N�Eİ �7�R���h@��`�(
��@�� Ё!ğ8��(	/�e$�A�]wb���?d)-g���#���(Dr�����C�G���!I�_��������{'{sK��.�f���P��z�>�7�Pz/x}�^�ʧ����f+%O)%�.V�>�9y 8�o�Y�ڢ�d4q}�o����V��؂g`�`࿘��u����_*�/M�ܛ�C�M��T��0=��������,�.^��_�������8&3E���1]����ߤaV*宣�K�W����?��P��|����������gi�j��fJeSk�$uQ��h�/ڳǠ��S���+M�x��}BM�9�+��rE�4dMӌ�����b�hp@���/fg�����Njy�|W"D��=P� �LC��˟@2b��+�U��=L;S[�1}?�	�c�'�z�ײn��Q��I�g���)�GD�!����3KWEc��Ǝ�YXG����w�W���qO�t���?�z,�����=#�Mp�����9Iq�����]fn�����\QQ8қU��X-�?�瞭���ܷ�Y�}x0���]���Y�c�����MY�W��Q����G�E\ж�aL��f�y(�3�_������ţ����6����)A�X�֕z�ΉJ+a��©�����\l���f:-��¹�/t ���'"�vy5��S��Y��u�èh�z��x�ۣ�ni{0xq�ʇ�|��_#[���%����*��5� ѬXX�'����K0y &�>�NTm��Q�׋E��j�@�	�����z�f7�*�������i�ǐ��	z�M��)+.���"}Ƙ�s��̥�b���93�R�R /�y5R��w�>�v������Fdt���v8���ډJ$J�ݜ��t�+�~�?<��la��綖Kц���x��+��0Z;H�fp�;����7.�c�sϋ����?L4j�ctҲՊB�뚚�&�n~��/H�X�A�uM�Y�����5�W���a奫�r��E��泑�'�'CR���:N^��#7�2�d&�o�ȩʓ��_���ne������;]V�	�%�R=r�G%N�UH	�|:��}�$�$SX9\:�H\�.)ah*-Ywkݸ��l7��TrCnElN9�����
��xwy�����=����$�a�V2?�I���)��5V��'<<'EI�I���%���-cO3:�u*b҈�Kl9�@V[�~%M���0`r�b$a�k�G�V����;-����m�'�{����6H��ca)��rw�p]�s'%���R�զ�ţ�L�L��Iծ���_�me$-:���y�'N|�ޔ /�B����(������\���y�I�f�f�~�ٸ�(ka��o�e�����{�)T�,K}!Q��`@6p���5A�`�҇��P_�3/A��8yZ,,,.1FF�Б}��'?�-_arFF��#��k\����~y�STf(JKI��efe�zQ<o��F8���>�!�lU�{�)�p�w���,.vj|?�!܉)_�1���ϼ��+{HQ�W�gmq��@WB�`aVN�)A,��<�:�^�Y��CJ,޸��o(ǜ ů��gwm�@���8Xt:U�.�3/_V�X@Bs���8�&�3�`^?�k�of�Z�0���%��2IL�P�������d�*�5�-M=���m�D��I@�)4�
�wQv".#(t"���k���R��,�WR�	 �ϓGEe%P=|��^;��_I+[kRk����J~��(�:I ����|8��d��%���z2=1�+�u���k!�p�P/>�/#�e�4�������5��D��t��*ɟ���8L�WD0�OD�(ɀ�6�a]V*�,_�r�קbC4�\ $�1�xJ,SR�r��z���oTgdS�[���C���m�:-���5�t��I
�KͿBʜ^%�*��'�����4f���Q(`���u
hR\.
���쳜��dMV�#�������IW=��x��1�ʐ�ߢ��3�����B�%L�D��!4�0+M��f�3���o��&x��-����Tl��d2��%E��`W걆���	�ε�O}�!9b��7���ʷ5���$˛j.�����K�8�j����#�psJ�{"��<|��[�v̆[�mIR+�?v��psL"��kDs�X��ݕ���)����2�_0E���c�3��Ȫ���ϧ����t;�	
�UUUlbb���n�F
66,�jA���IL]N���ē�E���((s�ak,)d o�~��oR��}�Ku=<��1��Y��t����K;y�V"(���n>��0��W+���,�P���sB.+ܚv�iND7J�M����w�r3����'{
���k�����-���4�j�cm\|\Ѿ�o�s(��+�cz;�7�������ⶳGԡ�5̙�~����@8�.c��m�� XE]m��� �0��a>�7}eY�՛ł'�äa�.<�L��ۄNm}.���0s������O�TUL��#�\�������.'z�	�:ڽa����H���x:N���w�ng�4���$�S����',x@���2m�]ەt�QO�ϧ��zkZ������ HS�f���`�eg_�;��l&F�� ��۪�� 0�A~�����{8ܙ%I�[��������灚��|��<��':�N��o��P�4L�Q�z�������4�c.�{6�?�2 ��U�Tv_�&y��v�G	?����W���4�apP;A��U�4�K$�ԧBG7�%[��r�6k�n4l4��i����=���d�0�����V���`���C��s)I�=�%/�4�u�9H���Q����'�,W��ЮY�B^ī܀��;��@��T烌(�7���v���98��Zݾ��1�����78HEC�xR�����J��	E'��=����Ϫ@*�^/+�:*��-�C������r�(�*�~3鄖>{�q�/���f�H�ܐyV]/�����ްd7��r�ߦ��0 �jfjn<:_���2CYV��Ç]V�v��+t��%s��k
/�w�{&[�s\4�)A�k�=�v���-7�#7DW�������"��yZ �2n����Ir_�ʗC��62B�̘�<�t~_�����Q�l$Ȏ����%>�=v��TpZDD���M�Y-�IF�/�pq�{Y���<���s�OW��Ef��iΉN���ߥH�:�0���(�8�n�5;�����;w�+�O�e:OG����\{�B��S��h8B�ޅK��NC?:=\K�{�����x�?#U9l|^}��r��'��c��)�=�Y��F"�쩅��h�n�x�ﱿ���ܼ��B��˧�pPx�����C�!��Gx��|�%���5Uq���pH��}*��^�{V��cq៞=����U>9��e�~�	��b�u2�++��pR�ȼ�굺�9J�ޞZdn��w��g�C����R�sB�x)�vb��/WS�֘Em?`�r,���]�<��C��H%�>�b��)�13tɰt�?}�2���x��iz��V;R}�s���7���&g?)�]�>^�>����c�����X6������I~�I�%���5EA�N���l�b���ͪ�\�N+>kr� 77���H=!��<���,�-0ߕ��D��II���"aK[|�|�3�e�_��z�;�hO���a[~���`�Lb��e6#H����M�M���*Hd��.^�$`�8�{=�r�w��K�~�y�b�x��>o\>l�{m�`/�y-w)�z)�ym����8I��N����[ �:x/�=<Ui~��.��*gM�E�77��El?x��{�&&nظ`X�iؠi��n_ن�8�p���n�t�Ab��K�Pd\;����.��o���BU� Y�%F��Bp&>�ß���]����k�k����ֵ�}�APy����5���K�M�K��k���r��jIy(C��EO��N�/��+��sU���ؔ�¸������Z�x�<A��u����d��:����t�`����zC�W��_e�.���������vY�S23cA�r����(hi�ظu��뒦/�T�չ�Z�M?ub�F�(n�f�-�u��>��f'L�������0��:����d����!�J"F����g��ɜǒ��9�*�a�2�F���������d||��>��hd����T��cw��J?~\�ή�Y��no�j2���dd`�n�>R~mH��D�ݦo�>?0�#�����c��E�jR��� X��<xkpE�fd��
��b=*�2 a�SW'@#��E�������|m��R~L.D��8��\��ݿ�Zj����'����ic�����'�B�5�% ����0���[�΅ʒ��Җ�3�I�R�R�_����)8��LLK�\����o�!�����~���x���C���?	E#z~��*�f�.ɫÕO*�q��ɡ�]4�+)j�n	�ܪ;/������g1e�I��Ӣ	@����n���v���}f!S��G,��"�\V�[��X�|
fa��"�L#K(i�X���|��S���r���^������G��R(���O���moMR��t�Z�8n>����U�!¯﹣�v7��76I���x�y_�B�������n���>?��|	J�+č��YSF!��8�|(��|f�C�V��d>�{�U�w(�xx�
�ď*�i��=Ճ���,��1B7�}|$������8%�A�G���j?�KȥBIy^���m�7�-.�(���EA3��3Ӭ��ot���m���Ә�N'&�2��ڣ�e~ge�'oY��/%���$t��j:�Y3ꉠ}�F��殺!��`��xg����ua6���T���w��j�2��KX�Rh8��2Yn�F�Ie8y��2_�&/))�R]�N,��M� *�� ���v{68?i=5�nD�2��ed�:�'3�h#"ƻpz�Bと}�R!&�����'4��[�oڮMJ�����������b��$?�_X�78���؋�U�D*�H$ǁ���I_�Dz�ɳ������]\\�L�z�����̒,eL�s���ꏈ�^K�G�L�?��.��a����贼�6��z�"��\�ęq^�_�*��q�h��{�c{����y�
q/mw���0��2w*�`��Ĕ�/ Q�4�����;M[
��L!X���kt��k��
�,	������D�qh�?4���r1�U<��֘썫�M��d�q`�+o�����4�3'^��S��$�vUGGG&9���Ե�`����_B`�����
�V��@C=��d@A�mk=�:i�ޙ���A%�oe���^�c��~_T}q$�B���".�g�de{��qX���.�􎏅{(~�<����r��ŢǴ�?L	��7��C�fo/,c��R���&kπw�o�ӿM[P߾Ϥ/���宥34N#�Me�O����l���O�MFe��z�Aڊ�G���p\H$��g ��4��[&�D���5)=�gRS3��}�
�f�fn�V�����T������bꞘX�.�g���^�����$2G;���M���
��`JJj3����2{QeU?�rS���fL�Z\�����tfV5��	�wk
"s�I��Ѳ#n2�_S&c;?0��{�6�}(��r�KZ���H�|;��& �����kdw�6��>�tC��-Kwк��R��˵���v�VzWhi�џ$^҉�	�:��l�s��am�ߞ��Cn4�	!�J]�����X�'Zī_��>�a�����zQª¸9�����B/n�Y^��.>��������4��� JBq���P9�W��+���'$�J�Z�T�L=�J�2B��B�x[7��_��/v�aTv~�K|闦k�g2��W���Z���صh�T�{m���:ָ=�/��W�%x�dP#G�d��(��4�K[�%���}�W�Tg.��� ��|<m�����P����"�y�9BIy1�s�g�Hv�v];,��n[���D��7X���?vi3��b��A����>_��9�ȸP�#�:8ty������/�+:�g^�~e'k�ħ"v���Z�����Z��{j�#���_���
�d�wJ�Q���N;�F*��*`S�"&��V����{�y��V�Hs�y�b�8\��~/7V���o*�֎j6v#g�{�#,�E�,��-��d�K7
�8nFA(�k�]%��TA������	����E�ʭ���Z��ʦi�D}/df��vB0RǮa�qw.�rx�pZݹbp`��<�Xx���I@�"W���b0;}�n��ZA䅤q���fM���~"onb�p�K���a��#����V�Ksj��l�Y�W�cBw���!ʋ6�\���3[��������|�}�ƃ[+)zP��,�UC�R�?9ϲ��=�g9�Rμ�|���@B>'ܚ�������EM��У���*���Gk��-�U��7��MwiF�K�����*,��ka` p\��;ط#n3�^�̗����D3/�%'�e����&�*�&�v=TWm��`���<_f�����֣L���fH*]u�%���tj��ҨԗRP����e&p;��p=A+V�2z�&��56���cf&xI��C�%?c�A�<N3�7�ԸEHij�R +��@s�)(`����,q.lؚ�E�*�۠��[����A@�����s;Rh ����d�x�g-mup��o��h�N8󜳿e-��~�pvlv�JL��aI�~��+aӿ(	3O�I�!3�,Q����#Qp1�;VW;4��}�(��O�Ϭ�z�/�,/O�|�i��%,���h��ƐF��>N��@8�C� �@+* #�\ ��sz�%����Ca?�����]���Ȫl�0�
M6�P��uϐRn�e�A'�W��B����څ�U� >�,䝚ʕ�=�	P�yO(h:?�]�\�@��zb����Se@Iy�y��yh%��SR���_:I=�(kl�Q���\8Ԅ~^�g씈�Q�v��_����AeL ���i|��d�c��ijfƣ"��/b���j�������(���{��q���Vl����FiG�&!��{��s���en�Տ)T���hZ;f�Z���ӵ�w��
	3�"*��l���22��)̫S�gѣi\s,��vAM��U#�r+r�,cT[e5�5��"��&����js)��ǓQk�Ro���h�6�>d�{d��T9�b�˒uڔ�1[���Qr��y�t|��e�3�5��l.����kA�޷{A�}W��}m7��}�;_�î�1PcE��.�k\0��Z�	+'h[�'��"w��O�^��3�#b&�t֗�Ǆ;&�*�H��'�]���i������K�C����umm'M �\�M�3.�%�G��2XΑ������H虙�d;`�[�Gq+�п'B�fk�p ,[�u��~PU�ɩ�ڍTc���eq�ys��9=n@����`�S� ��-ڎ͞�s|��9�)o�` 3X������ܺnG���;��RJ���ݧ��8���[;���+t�[�SR��)�������%w���ݜ,�=��@�����3�j���-�x��6�.8��4ᤎ%,�4f�=��30[�	�g*<?�����ɱ���UDw�Ɔ龠f��Rѹ!�Pg&�hg�����xFg���V75"�Y>�->���Ѧ\�ݑp�\�������Et�R�h"���:���3E�͑�ne��c�g���4�Au���˼,��-zc��429��/1"FA>���JX�����iX�n�]��g�����E�I�w����#"�?�yYY���t�H��u�K���sz@J����=�{Mm%~���lg��I��5݆�%Ɗ�0�3��FcI��1�`Y����Z����2��b��y'~;G�4I��[��eU������׎Z�G�*V\e�zM�s����^�!T�Y?��c����_q_���Z�) ��村���!?���w<���S��t��G�9�rc0s�$�5a�彐��|̯���?�vC������m�<��6v(��ZҐ�:��~K�����>�i�+�Ҿ"E!�$��Q��A���r�|����Ö��:��7��K�����Ճ�P�eWa?׽�u���Sޜ���bL����I�ZUL�y����\��e�۹�"�p��`���x�l�'�K�}!���Na�� x��Sn׋j����BQa�y��V��1_tbn;�A�l��z�����T�zM��0����¾^�2��B/M�8��7��f���n�h�m�tC��c:�L�.��͒��5�',���/w��}���%́�����MO�Kl&�œڬ� ���s���K��\Ee� �������+�k�RU1�A}y��~��M�O��:.h֡^l�!�����[���s}��/�Znv�vWܐ>�Z&{��.����)m�!���_��:�S+j���>���f*ii-<V�(Z�L>n$u�h`��5�A�GD1s�����z5�o��!C�����n��7'+�D0�\č�~�����$"tkpE���:�l��#e�w�p�is?��i(��a�?��8�%$З�%n���"�ܔ��Š�\Re&��Bj2�?���['2�\z��o_������P��t�}���#0�m����J}�"�_���c*ӦF���s�t�ڎ�=�.Ǳq1��KM`��j'��9�"��]E�J�迬��a���3[�ˆ���%�U8��|.B�
j�F폼�e��zk�(;����쪢"=e��BK�F�k)�������_	\c���B3�/·�bM�x��5mo{�_�b��KK�$��\�zHaT��& �P���9����Y�@�kZEE�	CT]?����u� �c"����������I�#`�U�Gd�R:םqm�z*�(��H��QaM�ڮ��2�r� �I>��;\����aGo��cf�d������l��t�k����!m�]3@���mM?U�DH��BF� 	7�wqOD���@�:�w1?��g<��;��%�㚰/�)D�*�#RI_�Fq�?lQN��T���,F�p%A�.l�
�~^á��j���gɵ_�q>���b�%8؝���@,*�H�
W���]]b�����3���Z�	=EK�"��9xk����ۖ�����r?�AYI	K]�3�g5W�F��Z�ZZ��gypE#��(!��=}(���gX~��&�/_�.)�N;ol�ޖ�رk9<��Q��4���N�	��Z���t>5��|�m�W�b!�`.g=3V
���3�z�c�_۽͈K�Zbw��2h�u�4�P��,�V�m��h����t�+]Б�K���� ��T3�|�_��������ݞ�> �$��3qm��-�p�~ 0���E8m%&/�C/4�uM�g��5ب7��=�ưZ�g\�Q��iV�٢E�im1
��NN_�}{��!��t�gy��j[5����v�E�X�ڲ���#��LH�*�zw�Iҕ����������$\�h�5Pn֔����%�E�ʢ~q��k�>ߒӠr/�	Cq�x�m�俙t�q>��M.�r���eu��LS�v/A\>j������2X&�����,{0dOy�#�oY��UJJ��-���q�{�F��CۤE�|YB�o����:�g8����������!�Y�>���c޺����_p0�0�B�0�� �H_.q�-��NP�qɾ��c�-��wD
6���.e����m�R"9aa�0�����IP�ԗB�|`�1��(��ZD�v�ߚ*�Z\>u�=ah�kq?]��'��=��&��Ňg�@�>Zح�JEl�,��@KK�*��h2�s�����eU��~�o{��e��ȭ������T��w�����qTjR#�7�$P	�b��{�dLwU��IS�ݵ:K�4{�D�l��?U�K��l���g��A1�a�D�RK�N�369��d��#9g,OΔ55�3�	;�j5�vmPa~����!���e�-�~l5���D �>6�r i��i���wY>y���ɍ�$��4S6�V�3i�&/I~��AT�_o=5�����1s��]����<��\�F;֖�V��ӵ��v��#7Ss����ZͲ����<Q��5XRUc���pRah�����T� ��KVI�]���'Y����U��+--r~�;t�}��' ΐ]ˊּ��f:���vQ�GWpskc�l֑���������h���/��$LH�C=� }a����Vg�⟕";��N�����J�z��UF&;{�DQY7�'���vЪ����YoƎ;%���[/���j�{\>}��¤�y�M`Ż�]<�"��**��03��ʚs �9ɕ����~�����(~��H7�LYƤ�a���G7ɽV>A���-��56U�K�Y�;��O~$�����d��c��y�'��0)�5�������z\jHr2%K���&?Q��wؽ��%�.�cN���~��s�ϐB�¹sPRWW_)�?�C�M-�z�����TGm��^욐�X�aŭc�F�(Z��O}xc�9����7h�Է��(���F�%��{y�����I�3߰��+l��]��Xܰ�+F���)����)`�Q�<hI��������Ia�S(�D6�c}Jl���O�I^�����1e��y�G?\]_��D�Tx�v�ȫ�Vѐq��>�N���C���mv�y��q�-���Y\BteU���^�=�L�{8�h|A����[�W�ݾ1����)H���r�m�NVr>%��Q�Chu�K�'�7�h~ˆ$�I��e���l���SD	I�Zs[Օ��ދDF%U]4=p/���	!yj�T�_��N��X���V5d�;��k2&	=<F��!����e\���>����z�$B�s&yL���P�$d�o"�K��%�-��D�a���p4�����''6�[�(>�W� /����m��7�_@��o V�R��>��Խ�,�2�9obleQEiU>)����qu�"0)�<��hΞ-�Č5N����V�Y�-ɟ��"&qtt,��|=���X�����-,�{1�����N�A�5��I�|���n]ƇD3;|Y��ޤ��Kᵚ-�ӷ�!�[���y��ɡ,s��	$m+QR)���i`K� c�:E�l�yuU�g���s��C:���R�3�=m!�r����ҥ�oS=�H. �N?�����_�%C��.�|u�:t�H����JD[],����r�z}�J��m{\�ޗ����lU,�m�h� �b)
���h�ؒ���L`lB
���W[GS.Δ�vB���m�<�����|v^��w�R�����֮۝��Yb+ ꀭ������*+SAN��Gb���z����f�V�M� v|�����*sj�Ȅ#mLJ�'�_>;/�KH���� ��_��:p�v� �R�xZ��6��Q�kL�f#I�3P�l���3?�qDޞAVJ5&�g�5b�����Bщ�]����c�aׇ�>��G��%���#	��Y���r�S)-kCp?�ra�ЖE�w5!u����C��y�C��|�5��71Ye#��=y��90�]��rk<:6��d�޼�QQQ��0̖Z��D�`�dH ߛ`<�;:򁚺a��H�]�j�W�ym�>zY��~�}$A��%�\�c�tDMj�\�*�oX��2f=V��tcE�ҘW��d�u�LF	,9�Y�@%SP��!ί�� �=��A��QP���[(�v��p|���R�m/��XN�")��`�+KN�j� <O�'�G�?�SSS?�Vh�6�j6#4�-��l7���C����hpQ��L��L����:�#��;�W�<�&x1��������ؘ��b<����3��z�zu�4Xe;n�m�Q�Ҵ�Ԩ����q���g��lN���t������1<����s��v3޵��-r���5�1���U/���D�D�!�,͸<˷��ɳݶF%Uվ.y&ʀoo����_1�ð~[M�����z�6���A��C�J���w7�ᱳ��~I�=���D�����!a���`�X�eP��Ю���z��tp���ſ��m�@��lQ�t��w���tw2���G͍��d{���p�H���5�H_o��uI��������~��qd�g�Z�\��N79�b���?��Qӌ1���ɔj�Z��2/�I�:�B�VE`
#���Ȯ��芰���]����b����Xma�U�گ	��~���e��	s�%�9�=��^�LT���}{5v	@kҾ弘�<K��<d)i�w�Z��~��2�떠�0EE.�k/�<(�Y'���2&1���w���eip8��k~�uz�DЌ����q��6���7�{X�5w��������=�`7+��"�;�K�F�;(�����!�׌�|/O��G��KR����-{�$�A����n/sɬ7 �T}��0S���,�;��h��rhx\x����[4J�D�糀
��R����j��g��k���F|��.�02��M����7���X�!��(˟_!m*������V���[��7����EN��0�}F��ӓ�v�z���vm/S�M�
`é��P����̯G�X�MfU}�苠�0���\�\~y�`k=#H�y��P�\�:��\aL�J��@�~�jȢ�\���^&��I��/ (�E.~���/����g���EU �z��A��\�(o�Ջe�iLo~C�bi�qq���d�f�H�E���Z�_~.U�!	�&���e>�2�@�_ױ�~��t�_au�	.�BE�N_��e�P���ey�;�6���|���8��'�`c�j�v����3�m��\�[e%[v:�D�M�5~8���X��~:�˙�ͦ�ذ��k���ډ��0��J����^�k�{���J{j�>�3w>:�|�9|��]F�ϭSE�'H��Ϥ;18Ȕ���o���X�ҹ�J��j��[�i�1�F�;31?��x��Gj��	qM����> ��v<8ތ:�A�b);��xq���ص/�5_*��>��&�����A�r1����[X4A���SV7ç�-�ȳ�Ê�N��6�������0F�N���'���Y*��*ZOX�F���7��Ⱥ�xV�����XK��xK]�{��z3+�P���{���Иl��Se0������!�� ��h�z��^x��4:�Iؠ�W��F������K��T/]��^��;.�i��}�"�'+�[E�1=UbS���ff�DF����IO�WUW7~y�լ6��͢�/�d��`;�[��Ubu[��]����JF~oII��D��[��w~�}���$~6�a`�������p����Ȃ��TP�3��s6Fntb]it��mѕ+?W'�O�q��d�w#��v�P��fD��5��V���U�jQ��Fb�Awe�����ȉ5��aY���Ԗ�x�\�M���,7Ϸ9���B]�O_�1�I�)������/���)��B-��������q���ME���~~0��D7�U��b ��gs{n_a�0���7u������-�%��t�ѳ��~�Qe��e��Df�aڻ!j��M��t�M�դ�̛!����[SS��XaTc��6�95H�]�E��;
���ȡ��e�����'�W��ĉ�����.�= m6^80G\\x4rbFJX7�Ka��2��?�lB��g�;�����CF2��f6o�l 2��?������O��C��ͷ�,��R�͘%��t>g �9��W%�����-~8����h��Q��Ͼ���_��:����iz\��i�$�)+X�-9y؉��z!��E�jV��$y[l��-���S3�`�%�wU�Ԯɂ�a{�!X��oap�9��t�T�]���`מd�$2��v�0���聕��b~�`��c�P�k	C�̤.+p���}*D(�`ؚ��R(z��0��h���O�����gE��*�s�_�z�Q�I�k��9bh�း�������y+*s��̭Y�wyP��S�N�J�����r�޵�4�,�3�qo�����Y��d�C���Z{۰�S|��+��ilT�4�)�o��m�>�sa
���{����d����M꤬��N��{��\7�g� }ot?Z;��X�53!wC��4G\�<߭��,��~KԴ��v��<Q�Ê��au��J�斈*�^�v�J�\	F�0�f`d�8��=e�a:{��E!v>����p��)�G��ѡ�'��ÊF��_X�޺�¨�v�@e T�)a�p]���	�!�ޘ�$�N���(ퟦ��J��wW�a=s�pQ..�_��hE�m$M
l��w���m��e�(Vo��S:�"��A�}KR��~��vq��t9.�31n�Dg&��X�p=Qà�����9r�щF�d3�IJ�k�Y�A�����'�G�!"��$�UX+��_����0-���:9�!ÙuQ.(�̺O��Q������t�UϪ�r�հ�a�7���/��d�4�>i��Ɛƭ�|ñ#��r�-��|<��ܦ�?_�>��]\�V�U�֎�+o�7��Џl&돨����V��|��R 4R�7���
��mA_P	�k���'��ǒ�N(1B'��.S!ɜ��؛����v��.��{�@�של�o�ݬJ�����'���%-�<k>DvAz��ZW������Emdј�����_7s�}�`.��O`��D��=g���0^����enZ�1T��RO|�R�������O�-����w��Z�^^���h $��P�`�0�#�`u�F~��>�)XIq���ѳ�W�\�Ez=9���}�Y�D��p��x����P����
�4b�z�Ί��><,�k%�xW(ˏ�+#n��= ��y�
{�N�|�}m�vBx0�j��3/��:���hxt�X�~;�	�&3�>s�_��7wh*(|��5��r\;c��;XS���YU���۠���Ki�HA��Ֆ�A�h�d,�
�Ǚⷂ����voW��""Bn�xbg=p\Z��
�[JJ
!��G|�aK���}�Uu�qy4]Hz_��x�TC!Y[oD�j.j�l���qz�Opy>^3�>P�b	X:�p����cll�JO��U\(ߋLKx��<մ���S4rn4555tfePB�*/��z���I(я��_�k,X��[?&ϗ�q��&a̫�ZM��w��P7��d�Օq�Ё��Ns�����;+�'��s�kk�OWjgϲ�������^Ū��9��T_�^k����jB�����p�<���[��܌a��ϟo_S5M-,�xx^��gZ	�g�+��\?Zݔ�=�!��{�/�oG�i��~B0&bc+J@�uu?�spL՟�w�׻�����C��~o��@���:��������u�j���Cs����#ŔC�AT~gg'��[+���y(��ƾKNM%�ۼ�HZZ:�ס���3:>[��ׯ6I�	II�;N�,gO�o^O���ޜV�Y�A8W.�VY�+�ܛj���R(������deŁ���p]��dU��]�G�$�F`�t��p�Bs�����k�7��J���\t��q��q�j�C�(k�E��m��3Z^���ˋ��R��!e�%�!hi�n-�y��Ã^x�f�U�p�И�ZB��QE���5�p ��bs��b������w�!x���z�� �db�0|���,���u��D�E�4ld'hi+���k������������mfq���:,�o�^��3��
<"s�yX����/1 ��ǐ�[��y5�P��*��bM��!�XF���9�����
*��Z8��Fip6�6�5��tMm���h��!͵e �G��|��e�!�]�)!�{�E�з�8Yi#fo_�l-�.���~6��G���z#� b�ye�DDN��_�{���_��>�8�zK�,�_��FH�����ɇ\���gV�|EG��<�1���Q	)��H�������v�ɿL�T����e���
���OG�TF*>?�g����=�u�^�+g�{��#����Ys^iRÈ��B����K�Ķ4��BeO}�4�a���y���n,��S����_!Q��
J����B���K:M�f�����]}V� �����.���kk�qg�͵�O;���D����
�4�]A@ HP�Hҫ� RC��(�{G�A��A�� -t��J w�����s����ݜ���}�=�<3����Бk��Ln�Zp=�.旐�/9�oڟ���ƶV����"���2�=��$ߧrNq�9���2w�|w��ר����T��&Ӷ��MR�G7g�{,���gl��W1�X���_%z�"�����-9�`����_^ِkf��;/�s���9B�^i2�,��&�m.��hN
y��2��ry��/��ƫb�L�����o�V.��ug5�"��x�y�m��N��'�)�)���-������az�H��}��Q�Ļr���3Z��̱�g0{��	��*�V�/�u*v�����1�|{�l1��.j�ɠ�.�[�1E��æ���(���$-����=ط����k,4i�||`��3Qi��s����師��B�S�Er&Q��d}rN��	���f@�g���@)[=�?�2�ݿ�&*���+�}��Y\\,"*��j-q��n�%&Ջt`-^��o��W ���7V��ƪ������۾�HZLѰ����B����QO����Se2��><�����h����&���������S��ތ5��Q��P���-�LHi�Q�]ޗ�WA&�3Q��Hr�U([+��<մeҷ����$;�k���X�ys�a�� �b�c�.-�Lh~tݟ�t��)y����]ccc7��c��5������F�P[����~T,k�:�mu�t������[y�|�O�l���]�*�/�b�$�(��Oi�`���q��'^�e��D�-��$�q���Qjt;����`�	�G�؇���s��8H�3aTI?q����`�39�����RBɝ�L�������x��l)���*k�V���ې�O�W��L�e��8�s�K�ɫ���@�S���-(���ȃ�h���O�e$ě%?u�1a��Sv�m�cwĚ��La��X�ZkV���s�p��T��93�::����w���'�m�ȴ�4�������kWW�t���t��'~k#��=��l�cv5���ו��MT���"Sp
QśUo���a��'1�O�=����{Qk���
����7��Y�zEE�~�7a��B�aޑ![gG̈́~Y\���pe,�d��w=F�+m9�l�Oj�3����4X�mxL9�	c�������r�^
��_
���.'�Z��8��������C]{�1�<���7�D������)�Ϋw4����d�,�f�/���씙���H�Iv:.����˟��Lyeanp�⹫���y��+���1�	��je�\}�bO]����g+��Q�Q������5u��b��d��=ςPp+|=v�;S�C9U}��TX�5ex�*kc�~S6Y������W}=��ӭ.eZ���&y�sx�0r���L:�/�(H��U�^+�-�t�h�Vii�?4��(K��>c��(W�����8�ZA:eE����-*.E���3�[�M�z�uk6��d=5��]w��xP{������|�P(�w�t��5twT@�����M9��n���&cuF���ju�Y��0�k�rnM���S>!-��;DF�.˺n��ڻ{�;�5�#����{�u'���S�j�����t"A)L�;��G@�t` ���hű��o���b)��Z��jas�����R�<���5Nt]M�c�y?N���d��2��a+��Ɉ�)�|+��)���ͩ��.���\��lD�Z�[�����'Jy�o�Ve�[[�U}Bm.ȮU��g�^�3�)�f�׈��,����������!�x��ֵ�Ͼ���1��l���P��lױ;>�٩@O�˯'/'.�S7s;%U��1�P��^��c�vD�񭣘��C�˃M�������]�k�,u�o
;aC.J��~<���zÕ���������h� .���(��,ش(zU;`�3J�ZI�U���e�ƴ���{�Q�ՐLk|+A{�C���k��h$=��p������@5��{�p�U�1Z^_�'����KH�k�^teY\�u��P���i�+��g�h�^G���UCT�J��/�k��y)��6�E�'<R�za	��������]T�|Rq�����1o�֑Z��Z��-���%e[)p��#"(����JJ�`�7�u����8F��hx�}{�Z��)9^�"}h�6>�$!+mo�Y8g��l9'&6��\�o,�H��6f�,<ג2S��=�7��!(��������b�T4t�p���޿�O�+y��gf�SU�2U)-�!�NҾF-%�{��2���w����U ��*��H���Zt�|o__�f�'�`ȳݰ�^�������ԴTۣR�m5#7���z�0c��E�8׳�5�ظB~���z\�b!�c�֙a�l�ܖu-6duoxh��d������}G�=7�5E���qs�=ѽ����$7���K������)��/1�,3{e���+�,IIIrb#�m�'%�������i���ui�[;/�Bo����`���ǿ�"�&��f�}��
V��]Z�^8��9|.�sĘ�ƾ�q������m��r��˨��g3���O�v�gEEE��KŚɥ��7=>�W��-J�Fvp<���4q��m�e�\�<:�����A����M>>��s?r���g�E������k��u���Wűz��L�����(��:vj�j��f}@ژ�ԝ�^�E��	:�כ�%&}��!�UUؒ-�ћz���������	�E�O���y�2�F�W�����~ȶؤK]437	����܉�8ڙa�a��p&RD������s«��r�e��1�e������	���Q�<�f*�^�$�S��RRپ>>\����/�/��T�j��+!�|�"����#*-(t�ǚ'��#L#�kx��ƒzx��E�l���z�o�"t�L0��x�gD�&�X#"�jVPPд%$�(�������r��֝�bQAal���/���B�_�6��YT�� ���@��+��
%�1Xz�Cj<׎�Q��R�1� I�e˼�F#�<F�Tvo��f�ƅ_��|���2�-�[C���:E�ׁ����{e�+'��-!�Zl����u���>D�3���P���>]/ 8?�u��7zЇBB��s)�*-!v����i�^:���MuJ{Y���]�"�����x~�4�Т��R'�R~9� ���{Ff�ERR��������?�l�I~}�޼��4�B�*9[�0V�z�U�/�<'�\~���,�R
V.N�|���W�R���ba$S.�|����S�._߲�ކ�s]3��w'+�+�����<h-�4��|��.��gW'��q�7�s�?�p�|4���]��*���2Շ�_K�f��Z���z��h�s뱝ݻ#B�㹕p���l��������1Ny/0G�Z�Nf-�+I��sj,��¥Ug�d�J�l?G�.����,?�wEi)PD�I��ܹ
��mw�v|Qt�y���s7/��0��}���N��«V���弪L\�nf.������o8�Ǔ3Sw�ϫaO������W���mgvTU{���vJ��/���Q�S�Ҫ�2��-_3W[�b����w��V���hu�x�hXr?5"�8pg.��[���e y*������\1�/�4��k%�/#��⾩��}��GĹ�L"��><�]������+��e� �i@
���:���b*��ꇨ���Gbn���(�A6Y��i|�bv���u����A\כ�����*&E���+�q�o��?��r�70h�K<Zl"�GW�KQ�oQ�:C��*Vڟ�1�l{ܰK�.�?#p1ƽɜt>�~�Х��N�&�m�ƮYK�c9'�}a�x�k�A�^'�����~�������.������*Hdff6��qRڇ�y��֛�`�	::��i�Z��m]���X��j����5��0k	��h��L�S�+3�K���n^`��L�7�t���A%l@k�k��V�n��OgZmA�C���l�Z�(�����ȕ�yߕ���α����C>��|����Ze���9�Sq�(��˩���k��P�R^����n��p�@Ս5���KUؙ���>9M���[[�����+@�I_�����w����0\�s��HW������G��G���kp� �'�ؿM^�h������H ����uʝkq�{"�56��$:KMW	]����!a�Ȇ��_G9,�������b�A��X-��=]]k����t���x{ץk�G�a�M�;��G���U�HO�����fC!���C3iǅ���xxy�^���m�A��ee�4M���Ȟ�nd4�m@~eP>h&���t���{K4��>�/t(?��ܽ>H�Lܛ�{}�`�Lf��뛎�<)lt���n��I���z\ߘn&R� ��ܡQ���{�@�b �|��÷�Rls��V]�����f4���
��T	���*���*vZJ��xLCN+|���o)�91��62� űKo�c�K8����W�����F�a�A�m�Ɇ[R�4�(휗+}2� �*��M^+��n9<˯��Vڗq�%_��y�uq݈K/F k�D�C֋����}%�xȒ���o���eGgqX��B���W����y��Oţ/�Z�g �އl��K@�&Ox������xT^ʗ+8^��������s��zc���X6�%���P�Z�	��Ǘ�\����@H?��g��\H��\��s���L������_by�����g��t-1R(Y����R�4�m�y;��8���㸼�V�����r=�v��TO)=���6�X��\��*x8���n�cd{�۸�O����9S�4��@!7H�MG����i>{�\vM���]���u�ܶ9�5E��jk{{��JN���Ae��)�fq�Z�x��[B	le���۸�IN=�+V��x!�CA�*ЦJ�w�{�6�s�w7�-��ͬ|�%	�VLMq��4�(j��U�1�95;�ۈtť��+C��E�'���/7���Y�y%�Z3n�c���:��
9���ٳ�T�j�q�h����}���r�ͣ�!1��d�����Z���8�?���%�4All[���
�=6�����W�8�}<��4��Y�φ��s�;2�یL򳒲��P���ɺi�_�.�3&~�g���>���4a�	��_΍�\����<�'%%e6ό07��ݽ1]8Z�O�T�`V��ds��Ƿ/�)����/(Z#�e�	�x1�����c�N��r�Of� vP&�&Y���r-�_y�Ʊ؄	*X5Fڰ���|D�$O?�΄0��b+%%�����R]Ĵ]�3�h�ƈU��I0#��{ǘ+������݄���o�Ĕ��l��M"i����ʼ�X����n��:H!(��|׸�B�a�Uj����&����N����[����AK4�\�f�_�#����S����;|��w)���+5�;2�<)��Zj�>����\8�F���������KVψ�
�N�*!]f��g�V8L��Vm�z�&�$N��Qg�-�A	)9���dN�Q�-�>	��S��g^�/[�r�sȋ���8��l7)�!�^|��� [��$�y.�CU�~��}�V|�Q@��!��xГ*�|g�ۂy�ש�~6daA�H(;ؕ3��W�Yf��+7;y.,�Ը82�S�>�z#_0ao���'�N�V�?PXd�&�S�;x9��i����m����m�HI��}�Q�_JI9@�+[��/bS鱕���O�KY�|0|n���W:�]ٵ&<L�����[#E-��3��ɋ��J�s�"�Bl�GӍ�_�����>�)�=��� �Ƙ����r�k�#Oó�KVX�B��.����>��I	�����X NQ����b
����
���ι�g��'��pn�.E��,���u�����-�ԍ6�]ʲ͆��/���Tn7ݑ�w�t�L����r_&������Sz4SR�ϟ��;:~����B����GS��S�z��?��oI4�m-�QLwA P�������*>��`Q���~ 
v��0�E��0�B�J(:��}󿛬����{�,��W�ڳ���0Y���p�������>��	tC򆤸����ԃR`i)���5II���AOP���������D������E 9�c �	���99�:�A
�f/����l�y�tt7U�=r���yz�����9ہ��X�����KJ~_�JdD�20{{���W�����o�玗��#������I)9�6� ���8���>0/89IU����� }����&��4�tU�Tl#�PK   �N�X��!O uq /   images/ca26ee1a-c8ec-49c9-93c2-f85ad300bf9b.pngԻy<��?�TN�r($t�Bv� -"KdߗL�]�1v9N%Y"[2c��F��`��c,��1�Ϙ�������y�x��5��뾖��܋w��/��v�����yM*��#�����W}|�r}������ǋ@���/��RQ�}#�?Qg��|�}��r���XR��pG;W��N.���2ר�nP)�?�v�_��GX�l���0?n~T��]��!gH�Jq.N����������� �ƍ�W���ޠ����dM�^O_E/�a�!<���	%������̓{2�]/�0?`�O����rgg�1��sZ)*ҏ�_Q�GO����Tg�G�T�Gb���=\���=z�h��h��3BeԤ���L#G|�N���MRJ�����H��Gcu.y�oT��2߲i�,�yϿ���©����-���7�r]�{"[��Z�|v�!ۣD��T3ەa_\� ���B��?����9%���KXxc����=
yя��?Î	��T�E����t�+F	|#K�h�ȧ$�oBo�<��G�:���}ޏ" ���R���X+��'�<�}�̲vy���j�MDx�J?-�V���e�^zJ�ڠv�-f���G\c����T�s�|^?+�7��6Xl+n��cc=���c���j4�Ӫ)�.7�����j̅�����|mzj�X![9���/�-�wx	��Ə��?�
W�~!�ݚ�~�Un7|��g8R��~^+��-£	�;��3�����z�K���j���y&l��(�Bّ�P΄��r�`�K^Ƹ���3y�������j��U������؊�ӡ���ʭ��\g���E�<'[�0)�N�ߌ1JqQd���*�uc���&�A��+�J8�	b��[��5�l���q�E�%dU�����Q����Ȯ��3#�S}�e�g����J�E�l�~�٢���,�$�(0���L�7�1�W,���1���վ�p����	)�E�x��;@���Y}!����ޣ!��f������0t1[#�!;�m���~?v���ǫ �c/�l���yh��0X�N��	s{)؃>����̽?��^��
�P����zo�����qv�Fފ\��o�H������� �?�"�王�zL'6�_2f�@����~	����W��a{�����
fg�ȋ����|�Id��w��DNtJ��`M� O;y�N 8l#ۈ9���;m&w���=q7�i0�v��������+�&F������p��V�}\(L���<ukD�~j����0��C�	(Ԭ�&1t	u`Ds���%����3;��[�ΰD�&)�߯K��t�4����fb9�ƀ�Uԃ���@�D��f��U ��_�ʸO���L@3�D�����.��,�k��2*x0��)���ݣ-`��l�}X�J�c�Xm��o��)���g�k^dd�}�pef}��e�&���|��hzݨ��E�nř�ƭm��o�\�	d]a+����[�� K�&Ʋ�����6���������^C��������n}��ƒ2MڌJ',�R�Ą�/ea�A��"��cy���kt<.\���X늟l^��B���у�Ș���9���@JX_�_�M6�w!�l����T3J̵����qJ�AP�m9�C�d��Ұ�����X4�ܒ�.��o%֣�**�B3ޗ�n�f/߯t��D�Jd�3�J7�/��$�ޤv��6 o��F�WV�`��z�sfUI�V'����7?45���3!:v�<Tc**�����O��A�GY�!�5<G)����M�#*ˢ�]S���E)�y�<����*(*� 7�m���.�ݎ���X8*"�����qQ�lm�2����sy$��Q���()��+]��9.��?*�,b$ȓ�%Ʊa��:6=@�!�7G���%'m���%��8G�^���d/��5���O��BoCa;h�E%ST;-��˱�{�{���NL�G%���(ꭰ���P�L9���Lϑ������G�V&	�^�'2�� >6�bY1O��ZL�\��
#-f��}xLh��۟I��֏���ۨZ���#U�.��;rk�o־L��!�c�r�x�Z�/�=���AA:U� �4eܓ�p?6W9��|֤���?�͎E�>稦&�0�xcA�����Zj&'kO���9e�e:Y|��a6@M��H�۩����9Y���� ��uA'�p�uG����I���������g�C%�z��Z�ϫA-0�~�8�R N�[�N�Z��^�M�e���i�v5�e�j��f��#5#��"`��ݔ\��#*��gL��) X�� �$����C���yņ��-�ͯMQ@�����]R3[�<\�v��s�X�<�����d# �k�7�����+�n��=�k�س��g�<���-
ﯕ*., e�ۣ)t`oh�R�T9����>U;Ae��<S�Q
*<Vh���[A�,�x�8����� �j��ok��;�h͊#d�/jzuL��U�������^|'�6
��i2�LFj&�%�ipʂ��@>md3#jj��I���h���}L��{��K�����n$�*JtskgN�q�x�u`�z�]n����%����O��DW�%5oX.�$���)|[;?9+@*1����
��z �
Y�`<^ XF��\�n�U)L���4c�$�5��H�1R�364�֘�NOl�I����L/�T�5pq&.GY{
*�g�Z�t�As�$O��;EΌ;?���T�,F��I�i��/v��&�4��)�s���f��JL�	�����Xو	�
f�����.u@�V���r^��G��#~�Ĝ�+6�E"�Y�V�X���̜�PR#�R��g��gZs@@W�^A`�l\�笣��*�"��w���s��3Ϸ l����|����r[X*����A4��Q��Q@�E�&堃�{�!�/�&�<�����q2؃�Deuv+ߠ�6�����u�2j�OA?��^��4w����A��v�9����	\N��'Ι��xo{��Lkq����R���P�2�|T_�B/�F2�������HЃ3.	Q�,�R#5iQ����N'��]�&ǳ@�2�?C����7��'�, G�T�{�M�yw�|��Yv�J��]M����n1ʰ 1X"�r�x*-�i6��f�6 � �5���T�Dk��{C\`�J?կ˔	�%%�����2S�*��h�����]E��Z
Q$���PҜ/���>�A��|:�F�P5�#\�e��>{��J1�@��6Bf�fy����� �yu�.4�7?<���>�z�S��hrB��̇�np��~W_� weya�
n�KZ�Du�[���P������*!h< 'c��e]������1���_l�����7A1t�\�c��K�IV5�q(���޻V9D>t�T+�dkj6�L���\�<�u�kG#J���yzO���݋׆�l�����m=>�)\���A�:�L���%� ��R������_��M�)��(�z�7���d�U��s�>�=X��޷�ž��:�s6�7.}��ȅ?�*O5��V �Q���p7�9-zhF	�<���06E��v~tt����&ޝ	,a��1���*p�j���|B�/�y׼l�p�	�t��Ǉ�n�%pg���Jb�+a����O'E�� �9�f��(�_�܄+B�o��9����A'i2K�=�g��Ś	H��+rҫ�� ��$��w��
tL���s��^����!���tǮѝ�3���s�?|����0��r��S$��2 0��|��1yoВ�b��cr͊7�6�8&Օ%�Ly�GP|uv0R˴h�.g��SzǸd�l[��2j.ޓs-+[t��a���6=!dwcj�J��X�U������9��EJ�@�s:Ȩʙ��&��{�C�d�Y̘�9?$.���c�a�����^��fL#Ovt`L�|t�y��
��ڄ��Opɲ�e������9$x��e�!��z�0����n����n�R�%��|��cċK�%_gb�ys���IŻ��g�Lmq^*�ѯ�����F.�X�z+8�	=�C���=fC�������e×���R� E�:��/"g)*�/׻���؝7��&|V.U��g4�� �ee�[}����L�9~���nܺ2�W����o9'�7��G8��+���P�␚<8ݸ�V�rp���sm\9���1�q���jr�4���v��w�>�$���O��}��E.��_�c/�5:�L22z���z�y��&���4&G�3M��P,/4:~+(f�����P�>	�P�����e6K�����B��j�q��ڮ���	��<��nX$���3�Ѓ��������
�=��z~�
+ל�U8�d�?��:a�UkEW�U�?B\���J0�a���������I��r�)m]����󗋧
���u��)��K�� �>07��	���uO�lG��O�T�733���*�T@�kQ@�uY4̅�5�h��]��Z6_ ���ȝ���=mP@F��`Ŷb=D.TLIF�wQOޫ(
m�hw5)Å`�7�\Z���*f����կ�t	NjQ�U�}�qh�G��d} ���+F���F�U��VQn�k������Ѽ�UP-
F?N���,zj��i��]-�t�7%r�s�)�����m�i"�MS���ܙ�>V,w�`]�r+:~��M��h]~�]~$�������t� C
�to�߀��+��-4o�`�c� �Fɒ��.�3qzj��؋�lv �!wL�XV�<Q�~_>�m���ɞ?���ש���@�?Rqn�[�s���;x֣8'1���Q��xl<��/�Y0���V��+��{�+e%�S9�����f ,wȂ���u��a�B_����Ѩh$ۤ���]`�>^�ŧۑ��Me.�l���R�I
�?lw{��T��W�����cR�޾����,�Y���>*�ls��]W$�������n���j�׷5�8�|���~7z9I�2�O�P������c��CBiB(Vsn3�3��Ҽڋ=+F�J#O�ȳY�aC��@��v� �k����	W�#�]kw^�����C_�űҭ����l����T[�Vfr&��v�4R-)�涖4%�${��4pg�s���)C�p��"�|R��+��'�L]�3���
���D]$ۄ��SIߪ����_V�]j"%Q�zs\h��w�1Yx�-����/�ڽWsgO�Bv+8�/�xsA~��^���{���n.��''�����-V�V����&o�+r�x���~�\�'��z���3�ÿ,u���x�^�N�+w��ؾ�V_WW8�0�c��d��RO�ݎ�u$cl����wO��6�Zo�x����1�!���4cG�ƭLSЫ-�Qt��[�y�o�CS��~AV���K1��R����{LG6/T����@���J6 �^�'9�	Y-�z�����e�C,����,�������^,J�Gm�贐ݘ�bs��Wk�I��[$$J�v��TU�/l���Hi���I�6�(�h3.Ơ��~����I�J'�d�����c��4Y�F^rh�oW��.�cY��6�t�V�˷3X��Q0N�YX"[�^�t�K�B��!|7K��vH����@餧��HV�5z��j�M��E���y�*����C�j5�64�&�9%/fF�p� ��8Zn���T���>
�4>���88@@j>=*r�Pϧ�b?݄��.jo4�0J,Qr�T$GB?q,�Yo�zf��g�X�|iV`h��ҧh���E"���s���6��c�c�3E):X �Tǈ��I���3������7-�נ[��	��I����|����H��	2�^�U.?, 0��ݧۊ��9n���T*�t�T\�� ��$�z�q**4	6m;��2^u������@��2��I��W3�'!OMl��Cqč?�ݏ��
HAq������q����Z���J2�l/ڥK�cm��Rd;�K�Y���X����]J���V�	x�S'5��N�<(��{���CO�����̙l�ި�=a+��:erMG�oI5���q�T�j2RQ��B�/�;t�E���^o��I��k{z�5B��ߦ)9��Y�w�v.l�| nďKz�������,��K�8�J�S?�2��\A���Aw��Z�#$߫3-�c�K���y��݊��v@���I��R=���;Wiޫp6MѲG�?Ic5�E8L5A�dD�Eeq���Cɛ �k����+H�X^��W'�`��O)����M`kM��5���60`0œi�l��K�����?>������-�1����j��s��#�W���{�
�YN�@�����7���� ������6��t��:G9t�3��?��)�j[������E��؏$3��1�ǯ�����b�n��Ӣ��nQ$AD�_������r�a�4�.*��cR	it���5�rJ,��+�W��1�Xs��|U:�|�7���3͐�<Cm�c]�
'R��ޱ��|^��Y�-�m[���w̝�\Z�pf�;�H��M>�5����]Jd����T���q'B&#2r\hT�;���"�?���{xaQ�^����\:����"���~�]���_�/��W�@��ܙ���Nw^��sD�'y�r��7�^�ջ3^m�n-�&J�%�J��h���PЭ)�fvQG�����i�����/��W���L���L>��t�z�> \4�aa�#O`	�
f�Sfur��k��cM�p3���b샥L (S��+Ւ3޾�0���M ������Q�e��Y����0>���\��a�9�x�?��S�ҵl�b��7Q��g�TD6`b�M�=Sy_S�U�2��6����f">��f���I�����Ҽ>�T(��C<9H�g);kWG׌N|?ܣ����)(�*��Ѽ?"r�i8��6@a_�)_�J��j��.�v��>�{PU�y����c�K��k��!Sg��W�8ʡ�k�v�OR����K�;ͯ7B}N���W�?�s\��(��8j��5��B�������@� ��$�Ks�N9��Um-��0���V��*��X�G�®�Z���}J��D笪֛���9�P��{�-��
���־0�m�k�Rl��2S�0t8ת�Dy ��n_��A�Ƕ��\zI�<`�b�����=Z�A�Nmn(V�ਞH��;���UyŴ�ޡo��4��U��_ա��wJM>E�oA��]��u�*B��M+���}��������S��As�������@	�c���=�TZ�s�ʉ��C����~=A��JRm]�[Y	|�Kgp���2Ӆ�X;O��ٻ@��/~�v_BȊ�����s��sXy�?&���d������y�a��r�8d��Mv=x�i���l�숅6;+�Ej�|�o�y��������'؏s'p�8�I�*�g1��	/�]�HYH����D�\f��y��|QL�,�W>�j�lR�x^:���%�|�ވo�8�h9H5���#=wF�o�Y(L��1�J5e��q���H�W���@9�d����C���ٯ��.nl"q*{N�Ro�([;TI����Vv�%�nX�ߥ�z�w�EV/G N��;C&U��'��Y	A��YU�+�سTO!}�c�~k=ɔç��>�A�} g����~68r����V� 8�=�j�w:�AGG-��ەU�Z�.J��,^W������|v��2=�K:cs]����}ik���2�gp8e��N%F&�<�;�5V�"&��I�u�����>c\1��ɕXZqA0y��M�H��4�_eE�+8W]��d�e�S6K�}��\�h���I�۲Hz��U���ʮ�����GgS����s��Wf��I9ڼ�=�t6�'���#��mƨ���h��/��a�@�����3�9H�����M��A� ����9^�1Rm����*'���	����M0�2N���2WN�3'���rY���� T̔c�u>3V�$h� `\k�^ۍ�r�0(.B�����~�(mR�p)F`�+E��	�z�p^��l�r���{x��*/\��K�t�����?d:H����э��C����G���eW=�Q����H�P'/-\�39��=[�w��]�^��(PQ�'}J��
L��������LY�ϰ��Uo7΂Ճ��}uA�1����}�:�6�C����MM��z1m��� B�|?啒�&֔r��<O+�C��ܓ!�'R���S���g/��_��)g�¤����Pk92����TKd��}�bM��?'ZA]DCz��j�Xr|�y��5�˧Q�V��5�r��UN���Dn��E� �#��Iϔ�fM�3�xς�L�M�v!=����<K�CGz���/�3��¤g
��3b�pl�������̣'��?�9�.�Q��
J���*6����q:�@i�*�����Nj��fB8��W1��#E�NX�>O��8�7t�Q��Dj�x������?cN�(G=�(jk�.�=�W$���u~��_fq�wp���6�j�n2��,�����I��o'�2��I!�a2;�N9���5���@�Ao����]�����i�f(�J��*r݉\,�͍���� �����-�p��)l�Jԙ��K�l.=�C��1`�z	�u"���nL`�{qbQU��pvm���J�q���KXR�$��k�um_��Xl�S�&t���!T���ٻO�J�r�-ڲ����-�XJ^����#��G�#1L�s�[���fJ�54��l����"Ɇ��։�,�(QFQ�e`�i�����VA|R��� D�r�D&�ѪoJ P+��KS
�������[�X�����Xn`�\�E-(a�
$8B�!�_O0PF�ٿv8�۸=<��6���)�4��2���cR@nh_�4���.L޶���#w���| �Vǁ4=��w�(v`�r.�+�.j���"5��;��9��^;9�>e�O�N�lV&�4E
0#�Ɖ�F>>���V�ǎY��T�Θ���2 �1���L����e!Y�vDl��`,sJHp}�w.���L��y�n�ͰD����h,�t�f�S��<�hc���)Ҫ�6y�`�>N<F�ٲ)�=����+@DN�;�)�E塡�軼a�/p
��j��@�e�'�3�<x�����E�t7)��1��D�9&,T���ˈз[�S�S�F�[1�^+tԐ�+�f�@��-Fv�)6u�Hw��n�ï���5F����$�
pk�ŧ��~y(,
�z�r�Q:�����N  Q6��˵]GCʜ��I	>�+��<�J9����j؝-�n�DM(0w�o~��|C��W#���U�af�3��\�piS��\�+�h�r�J�PY;d8�L�Mq�].�9�Dv�Ro4�%�\!n�Ƒ�L���?�B#�_��1�M�T ��(��Vз��V�������Jh��:�a�w+��#�!�-c��B��J1P���Q�g��3���&厡D��X�r���J(BX�m��:��XU9�5�\5��<{;o�t��"��٨U��ى�ЖH���Ԟ�[��,��^��LKxߠ5`��ȷ1�?b}��L�*|nrt_*XdcW�~".K��C��"��G;C�c�-eo�N9&Xs�������"�A��"@ Ma�.�����h��]���/��7SS#��(WR߈V�M/x��)nG���j�����Ub�e�\�hd�ꌻ0����z�0��K^��0�]���U������,��	���=s���C�C3~t���#v�����,�c�ac�s�*:�7y�
} ���c��ӯĆ�'> GG�����k�.+��
�X	 .����R�fډ��`�����`��K�$�dZɇY��*����C	� �<A�	�8>�}��`/Bx�t/f>d��9G�vU%�������MYZ%�ْR3R�(a38�c��Wx�w�N�YP�n�����������r���#Y%|�ܼ'���Oɉ�6�.Jt���W�Q5~�7����Z�K�p@�W{���H�8�n�+��O� AD-@�=[I\�a!]1eb@`�d�3t�S����a�ؤ�t�k:��̗>���1�G��m��
e�DV���Vtx�\k�Fl�o�������J����q!�`��?0��*J�=v�%7��}W�FN�I<b�"Q�x*m�2�P�k����F��ٍ���>X�\i��G�Xa%�d����GS(���Z���r79�:�5qT@���_A��M6E)źv�)l~h"q��,�Et.j���Um�H�H��5*1{0��h�ǝ!�Si_�X�$�c���]�kb�÷�/IA[�H�ȰgUqJ�UB��!
�gI��1ʞ�c��ّ_�i���I�&n��HJ;>ߧTbĸ��b��"h��r�������l�J�|\ �D��nm���|-��i9е��p�G��r���ƞ���xi�]sM�3 n��4ʶ}k���Ktt�5�G{,��jV�z�C��� dNP&R+�r�Gg>��s[��q)��g��ɉ|˟��*�E�9��Vf{i X�(`�����(1�c:\�S�����ܾ{���I\��iE:TA�\GR:���f礧&%����H̫�F��_h�.x<X��IE1�ɛ���@Dsr�.����-:��D?G���g����T��-\��/���/��|zF��Ko>�j����[�g]�/.^.9��p��^!�X^�Hg���D�dtŨ4!��e�]��?ٸ^Q*�׮�^$��µf���h�1R�����1� ʂ�j��	c�W��u����tJ��&���M�b���=���	S��^9~T{ᷝ����ԁ��!���{=�(��0%��G9�r�ѷ��x�)K�N�5[{�X�-¯v楪�����*ß}}<�sg.i6���t��Q��K*�i㱐���_1T�*_�����M��)�����~�U�)��M9���V�����l�)A����-PT�/�(���}̲�����������=oQU���^m�{�������6@;`M쭳ETv���=B������lߎm  ���/+��pI��%5��E0��\�G86�&znO�Q�U<�s�HumIm�3��$ÔJ�X⢏i����3��"yyE�H>A=� |L" �0e�������Uq���À�W.���/Gg�U�]�l�PI:����{7pYӗ��-&OE	V<U���r	=V��u>k`͏���;<��n!���֒�!d��ONE��� �U�Xg�����fL��}���u�mڦ�Y��О�9�W �5Z�Ɠ&�|�A��c'��;������w�R\1����acR}\R�M����Z�u�ҋ����G`�>�晥֧���2i<&㴰��HNy�.j�����g���NM��zu���^�ιR�υ�?���k�f���쎭����v#���mŚ�.5M6 �x��֕XA.�>��w�>��ޖm�3kg��+��h�T`T�~��W��ϘHFk�A[!�������K1���3~ e�+1;�<6Y�ٳՙ���P	���ͷ�=[�}�W5K��͹��ˏc����U[��b������Q�<�}��on����	,M��{X�?�l&�7X�U�ά��Ϭ���#��IDf{�GO�����2@���l��;J�MB�  ��y5.lF�Yh I���?2{mk�@��̭M"[�_�W$���n����<�5V�0��z��#����%�P�aAߌ��R#�S�>�&X�qg�X�����	��C����l ��c'J5�Q���K�>��J(��"��^�lM��C�I* P�L�§+|9*�^^�Ք�sg.|U���R]6�r�&!�$�+�Î@���E��2`�(�t�: �f�K� R��h!�Zx>�����|Zz9����K1�|5���ҷ2��}́A�ze�'=��Ye[h�pɩ"�|� �Q�VVrY�P�����Q9Bo�aË�\���!����i��Ľ��W��=��p��hA�]��]���ɢ���+�B�z���4|*=�9A��r+��8&�Gwm�l[�[D���ʝ�+
2$��?~�����6�FU�����3Wp�lw��y�����{X�9Xֲ�������n�83%�T�fv��r�ř$SS������d���3�S���n�%�d��� �^Ш��쨹bҞ9қ���祖��'r�F����%�)Ɉ��7V�ӊW�b�^�^���Ѿ5���8mz��������p��*�Z��m���0j��Tf�4P%��Y��UqS���'� �����jt�����B��-���/1��{��liY��L�XA����}7�K�	��Z]��8#�tF�a�s�ɟ�d`]>qaY�B�t(5Xzl�U���|�j���l�F�u�fVޙ�^w�)�(�Es�5D�D"un�qԥC�wJ�9Z��Q�I��^��&�-d�H�,�9����W���Ґcsq�H�Zb�k�XZ;b��,��[��n���������������x0k:?����~�v�,1^��fuz+����{�^�ܹ�՞��Ő�0y@EW;Z'T6u�i���W^�[0������A2�։��)�;��lz�4�JP+2I.1�=ã.����79������@�p[���!�9�uBz��������7�RaT�u���:g���Ů!x���cA|��WϨI7�v��S�d!�����	��Ͳ'>�5��w�0_?*bZ���9
Py*��)!���jB%MFL�����Y� 8�n>	�8R��v���(�9�<�톇�t����-�T J�F�/ _��琐e�X�=C���	�(V���	��6�H[�9y��~k,T�f�x���1�i�&B���eh��؍�pm�hخD`0rK�y��"v<��X0�.������#�qs���L�S�r�O���jF�5�arn����MF�xǛ`��,�!�/�H�%��*�d;�����Z���Y,b���U�:�.�-��Kd���$����eإ��Ξ��
~�M�?������_W�aX-����^P�Q-p^����)��	�`���%���,i�E��_<��(䖭Vx����Lf;���8��bD� r
��Ѕ����e����y�6�<ne���e�%��@��0��ݐs�;AM�-@���0�@Y�����%shDJ�Fk�GhR��4�^M�c-v�����������޻�}\��Ws��ݜ�L�6��TV��F��J����n���:�S^��m�]��'Ο{��FI���\Y���:^|c�b�F��ss��$�Ձ������_�ͅJ������o������3��O�uv�h�r��7tg�؟	��
S���j���r��gs$��t�&������"p�i����kṕ5��e��>�вy��̥�V�:lTփN�%�t�3�؏�|��� /F��`�1�e��s�¾C����^e��Ol�f�q�kJ/>WO A��
��=H�Ȇ8>8��!��S1�k�:���S��)N���i����L�촋l���0����E����ٟm���y��X��B#�=���j�zG�Ƿ��mD�*/1����y�ç�Q��2W�@W��%/ޚ|D�Q�_7�`�m����18��u�NK���Z��Eپ_=���d�ң�-"j���ԑ��@X��t�p]�	�O���~8t��J����ڈwdkX���w�Pz��� jx`/V���32 �&G�CznhAl�����(!��+�=_*P���q��ʗ��ǿ;kN�ӕ=��c����U?%3�_���)�iO,W��I��:�K���T:�6��^l�|J�wa�/:��|���{6���ݽ��"���Lk=���
������@��<�F�X��!����ȅ|�x�hݾ!��`X<9�m�g�v��#���[�_§4+LQ���?Ιݜ.�^F��:_��nu�e�J8�Ω�&j�������@P�jX��o����6	u.՞��ߌj�:��}�4��0Dn	��p2�$�Ql����tt�%-�l?��p�>����q���oСT+��n�sP� CtE��bD�LC�vZn��'Lh���|�r�i��H��Gu��*��U �%l��-G44��i��C�A^���>��۫������rQݶ���c�v&.�� ��� Ձ���p���Kj�3�J��[��?���A�`Sϕ�5ӬJ'{m�7�)nZ���K�l��������W�ŻPT���J���9���3:�����nt@�����Ҽ�������k�`U&I��AwU�'c��g��o6�,������8)Mn0�X�;Q��ݠ��WքE�OM�m���hQ�q��E���-*lo������u����4�g�盚� �u`� -0xi�fa�R⟕]�Kt`O���3�H�����q���"m��m��	�𻀍��[Mˏ3i��b���c��64��u�jV/iSDo��Il��Tn/�*��D�=�f�$x	=�}\�G��J~}𷶒�f�YC��'�7����R�Mĺ@��@4���~ǫ�/�,����Ë�~��f� z�*�!�{��D�!�voc�ayȲ��6ć�s{L�JF���ssĉi��jg�Ҫ���2ˬ89���uf
�5�/r�5^�f@V��>��<���Oj�"��Po�3!�ǁ��Я��\=#�xK�����"���R:�>m�Z�Yt��ƻ��Z���3ĺ����j�4'��&ޛ9y��I�� ��^k�b��,gW�>Y�Aiw���}5���R'�nt0  �(ZL~7$+c
Q���j�"ʴrB\]D[+�R�^��\�v�o��!���+�3G	;s�(K�%�f�E�{�YU?�@��|Z��0GuȻ���3g��@E�����|öz	��b�������U`AQ��"}��l�W�v+Q؈�1�j�ի�>��N�D2T�Î]�x=.��c�)��r�ʫ��FJUU�@�+�wi�}	"��M�b��aJ�ilEt}���7J�aI��m�2] ���y�bOu,����G*��<|����(m��Qy�������C��oD�J����#N0Tžxrd����G�+4�O��qb�i�)ń3+[�#���%�����p�t��*W�=���ۓ�(��}�'���K3����E��++�֟�E��TTck�i�Tؙ����s,���^K��[�+C���C���G�;y�j�kj:k�����%
V3RĽh7G�����T9:߳O��hS�Х-�{-�H7�W��A����W�����2�g�U�zl}�~�Z�MDj�@?'�{���dv��}R��+�����Y�yK1�fb�y���̧�?}-[z�����|N!�I��������h�Ѳ�7_䆥��L�Zl�ᰉ�Ev�/�!Ϫ���i�T�0�zJ�?�� ���R	�V��/�Z�����_����Å����� K|<��pg-���MIe� fdbb"Tf���g�pI0|�`R6��TΫ�M�ȗ������h�絎�����NyNd���+�:�����:"�f?~�hnE�a��?��:�v���i�{2���c|���*�Lc��4�i0��3���mlRh�S��&j���*VrO�����0>�X��������_����g��Gɟ�{�e3�m"�Jr'(�;!O���r�v��ه�}����;��g��¢��j���j����޵j�����U��T��m.��!㽞�^�;���r���7q_*g��}vK��U����Sc#r�y�P�I��S�ð9!�����	���a���@����~����0Ot�Z�2��y>zE"/QڴN�Q��n�p��7|�;���P=`	SXtϣ1aR������Z����?&��y>��\Z+N�Oֹ{��	)��J8����7H�����o?�1�L�=�Q��z!c� ���\{M3O�S�>�L���� �8ZT��YJ��(����p�����]����O��6�#v�{t-�kŖk��(=��3!�S�g�>f��4H��� R�����g�����X�)�`��O���f���>�q�lE��6�ӑ�w�7<��'(�.���N�^J&`�񹟪'������{S>�eb*������:��t��B�.B\u�S� j<H���m��yѵ8WOnf�4ђ����}�byq}���u��m�������Z5N1���8�,�Gګi$��Y��!����= Ƽ�o�-�(�{i�a�3a.B=O�3�0$bS���S�Q�{B��S�k���i���������կ%��g�����G�5�/3�K��me�Y
tڈ��ya��@Ԏ�^�Q����h����q����k�~����]�"�:̙iU���=�ko�"<[�V��M��k<[��PП}̲�w�G	=?�]+VWiJ|�9��NE�</
�F���͸ql�ho, ��Zo� ��.Qu�^j�绌)�ݘO�'�o�| �i����L��Mۯ�"d��k�]��C|l>��i��`���!����@���ژ����C����4+Ҏ��?�-z�9AEU�[�?�]�Ϙ�g�Ê��n �kW�>�vzk��q��~��/hq
J��h�w�c����/Xuk4��c��e���>)r�Sg���L�&��o�}̒n~X���@�[�"?*����m���ilЕܱ� 8�bD��4�y�)S�q��1~��	>��QTI{�#ˆ>���i_���5<틎m[�.���|���W��L!�����,�`{�����ICO��9�ߋ:��/I�_����k���7Mh=�B�?�E Ĳw�q��U�Q͍�]<O������MLE[<�GZ�{h?�2���T���/'}\%F�1�S�K]%���"#��%�$�a
������ 诂���O�����/��"6W:��{�O�	��PP�M��_�}����]���=X�^�Gڏ�=�T��22�
�:.�� ��	S/@�rOv�;bW�C��������M"L�g��v��h:4)���������kO��Y~_�}��Ǫ����>�KZN��כ�|L �-9�0�K��m��Ѕˁq�"1#�%��!����	���)�_�N�T/��׌;�Nܒh����s��jʊ�������x�r^8����V�x���K({8�>G��]|m�-ݹ���Xj�z0�Z�3(�W�8��:"�y���Oj"�i����C��]�
Q �Q4R��|��B�����v��E�̊/�T89�,�֬��3_za�$� ��=|��|�yt$��+ e�@z<�g=���#p�1�o ��2�^�/s������U�[V�?Ύ��|��K�;Ab�7�-qɩ[�������l`K߁�C�^�UwS2�;�t�1pe��{&hR�f߽� ���Cb4�Tr��C�P�t��[���p��m���єD�eq��p�܁P��ki)���(�**	gWE�8�$��lmٛ�#g�����wٙ��eo�{_}����{����|^�#���?%)du��B6<�X�SK��L�%QY���
�'�|k����ķJ<�_��H�{�P��o·�z 3�l��Ԧ�\U��<d/��;V ��<������H-��PP���*�ɫP�_�WlA�BW>ٹ����=6t�$�$��ɰ�WD��0�I����_��������[�x�ZG����.�}ٟ���
�dvc9�p]��ߩ6�ՕFq��������A���j��?���)�_��*O��A_9^�%Z�6�uE8Ȣ�k)�<iQMg��� �N�̊~��^��n?d�wK��%�f;��xx)���7���j�U���Т��	�"e7,�Z��
*�Tü���D��
�:I56�s�:������O���l�/�4�P5�3t�-�{zQ�c���`�;�l�'��n3�]t(� ����\츈cm0��`	�ޝ�ju�^�+�W�E�/�i��.�B�8h��rU���/���S'8ޖzL��ÿ��>�&�W�ɼcܹ��������z���ǧ2�H/�Y3����)��؛ǔ��o1�d�DN"���)!�2� T%K��Ce�q��M�Bq��Ys壘ݯ��W�J�)�qSS�44��Soݧ���5>mgW����Qop���°!t��������
j�i��O;��-�J���v>�|"�6��cZ̢���\_�K�6;�bP���{zV�V�� EF���䣩L��8�?\}�δױ�d_�f�0?)�SN� @���3���=)sm��d�Y��.���}l�F �w�d�����k|'���� �Z��Lgj8: E<X��#nD@��-r�����7���5k��9�m�0�u� ?�������8�`/���_�6�;���ئ{-���y `�pf�����sCޓ�b��ʿ`������a�ڰ�C�y�������*�8u}��=,�p�Г]c]�a����&W�g��Djq����,μ��f�;-|<����Jƃ5��E��}�R/�(7�z�kt(��k-�ǯ^��/Θ#�-w�ǯ-��M=���3�+ �>"����G�>a&���4��e`i����1��B�QK�_���$E.����9>��˱vM��#�>|��[���N�-�:��W�H��ԂA�M������7��0?�;~���4��p��7��� �>�u��ep��(�~x���̾��a�{�#�����CV~�OkJ��J1֏����Yv�z�(I�����ͧ�@YSj|}wwu�XG��%E��lr¯��u�W@������boH�t.?l��"/�o�����s���0\	�z��n��}�kнBEיr���'OAl�����+��ÙX�7+p==99��ֆ��6����}��k���gi�	w�Λ��Rw�<v,%<�쁉NG�_���v�M��
A@]�-E������w������bЅ������y��a�$7�������lU�5�i���ln<��4H���Ɯ�f�gk��K�̃�,h2\`i�p	KkFs�xw���)R�<���ުź�Jp]�O�R۟`�C�(��^2��C��`�����,����������m+�.�8��������Rc�� G~h�������s�(��e�|�%HAut��2�===\��,� ���,��=[l��E|��|'�m^�y�����fv�%�oy\ l���E�a�R�¨�bؒ#�!����.�}�t4�3���G��z�
�0�����q��`��ex�Ðʻ���0�����4�/���pn�ҭ�5<�IU����|췿ut]�Z�݂�-�OI���Ш|�� �V?Q#�=Gl���s������g����٘0��ׂcy��:1uoq�j����l��Sk�pl�d#f�=a��b��@J�*��<3 ����Aڬa�).�_0�����{.�~���'#���tY;���+v�f�[W�r���7���s�2�<�uG݋F������F�*�8T�bp����DЇ�W\��2���	�7�A`�|�8U�������B�+���o">�ʒ�ULP�*)��D�>E�E�)kt��}�������`�%XOr)�������
���m����a O1������=�q<���e���_O���E��v�����,M���|5�x�9ތ�ve^�h�����h���0f��'�II`�NO��Z7�ɯ��qy�LGr�F�q� �RL��S���<����`����_�`�S{.[eJ�fiO2�y��mܭ�A�%]A��?��4%8>��;���@�t0�.|p��:�<�����ߏ�.�������u�n��H"Zh<�m��CaA�]�qa���h��g�����RG�9��t�V�N��+�t?�Ϻ��_�3�R�z�s���.$2�P#�_R���(.����ⴙ'b�,��u��Q�=��K��u~EO��e��!$�;�F�L�lrT>bx�=�3��3~�{!���)���;a*����7��U�N�}�?��u��ёIxu0���w�[�2�Uކ�jR������v�qP;ȝr�e���]72��� �18��Ϯ��l5x�e��	]�� /��X����m����#�iQg��k��g��]��kɈ�e	l��C�M���e�d�2=������[rܞ�Nv��|��-z}�efPe�l>6f�[2�pV�Q4�v���K���4��\�)��?gh#�����I�z�Y��C�z�_/����쥹u�'\@�HZ�n��%��o�#��
i�.���̄�8�N'AC�*��miV����d�u>�GP�q&®����P��;�`�ҥRB��6�\��%1��0U����3=��'?%�}��[ua��\���ry
����藺�y�=�U�u�ƿ��Sϕ4Et���䬫,��e�d�~�<T�+m�S@A�5�n�ӝ���
���2�����C�d
˖�]�E��3�w3]������M{m�|Hx�b��g�Ã�+
�����A�C��6?�����/8X��9_��Y >wZ��K��:���4������B��}1'��eS�m������tgd�z���,~�o��	S��Pn�0���*���U�<�/*l�7~��.c�
;1�����dCOd���lg߿U��(Z�h���6�G.RZ!�N��r.Z�t��MpR�d��k�ؘ)���Z���0&��=�O��n}ͱ�
ެ[�8Q��瑬<�~.jB��k�6��7NS�i���ɓӥĞ��VL7�*{w[�g�I��X�H�~�KSG����F�	zZ7�"�~h��Mb�ϗe�����m�3�0���1�s��3�Qkы���ɝ򑷋��?Q��W���Y���))�3"�	R� �a�+Zcţ���W78��G��y!�w\�T�|Б�U*O>�@���D�]��e4��h�u�;�UX�/%��F&ȍ��A���ܒ9�r>��i��E!S�$X�|z��i~���E��7,��4��}���*�444tx1l����x��V4�[:Ts۹�1��j(^}�X�ٜ:&��х�xڦLP��N���e��,��J���u�#���n�.�G2�vXO,�d=�K䟸�k[	����/Y�-����x�?��$(N�4 ��9&��9�A|q��|�$��ڐ�@�]��rt�S������QB���R�
��tx�}�cs�-�|0@�Ε[r4��Y�Pz2%4�c(�UxB��p4I�l���2+)���]���T%�I��1��8�f��j�N*wJY��}1,YJ$�%��%��t�?\v#13��8����7'Y���cm��`*Z�����,w������<Rc��h~��O[����EL���gG���y|[��t��І�Ԙ��;(ɯ���^�y��`\o?�à�c���521�ɼ[�ߒ��<M��b����A����ː�,JK
�K�5I˓GHR#�]Y��w�b�Ü�q"%�8y����jć��J*Z��a�Ɲ��҇��}�t��wF]��1��"�x���|�\���Ϋ��RM�C���_*O7���Z�Zmw���j�`��x}������v�%����Y�7�@�?>u�L!��T^���q&v-f�tB)I�
6�7�d���x��ѾA��BN�,�C8�z��"�t��'���m��D7K4L��{� q�Ұ���W	�!�B�y%�?¤];tu2��q����1�r�@���gY��8:2?X*,}���"Bu��Av���r|�֯��+�䐻�Z��+�ʅ�Y��TMwرS�c���Qv�"A���ǷR�=�A�!wlK��ʯ��:��u&��PN��p��[��>������[�'o)]qЬ�g]�g��L�C�t�_�5^�+Yf���h˸m�dD��p��H�7�A�t�<4-4]�����1P$_�b��w��V��hq���O��E_ZjI1�{hײ�|��R�&��ʧ�ް��L��F�'B5�ע-ʷ~0i:�� �"�K��)�z��1J4YdP���9B�pf����}�)b�8���������U�|�F����Z#Îς,�n��.MTCJ�`	��̯�����[Z6�v�0F�o~�"���3H�����9��K��x����ş|'a
e%h�V��(o[��5���;I/���d?C�hCD ���G�B�b����QBCԼ%��x]R�qd÷b?�F餩+/V��� �ǩ�Js���a�H����}(�� �U�
{!>�Բl{x��� ����'���8������]$Nݙ�W�ҔeK����<-�=%V�-�b��(��J�X}��f�v\�Cd$�W��
�/T�v׫s��s�?�|'O��^Ei�����0�+3��
���"Q�8p(���P�D�S�#�����}w�g����Mfk�d��&�y�$v��bE�����D�� Q��gJô��SP����pJ�w޵���o��%K);�=���u"�.WE4����s ����h�Wl"��(}�Kn֪cRs]�Cb�TĮ�mb��K3����:5�Ņ[���
:/:��Pʯ؄FzW �F�KⅥR�Z���%�g��T��.wXjEoc�91 �o|���t���4c�����:׬�����z=�ӣ�	������;1��`�������w�Sf<��'�E+"^�?���crz ��d��!�_�Ѭd�R��{_�t�nf�<C8h��H)�r�3Q�@c,ʇ�h��6�% @)�-LD���>�z�Cu��~l�%2��=���)d[�SUرv3�-���x��(O�aT�C�R��#b 
�^|�������oU+��ޮ�����y\��v,������Qv��E��%��ac�{|F4L	G%�õ��û#�(���0L�JĲ�Q�UyD��d?���A��R�M9�o�ݏ�JW�����B���Ra9�S流j��;l0%���!����� \�ʕLb����Ϳ+�,.gF^�R�s���Yvb�_۾��U�p;�\��K�?],����n{��Ί��؞VM]g/�6�2�m�T�q�Z�TU�����8���t��H�e�ǸTŵ̌��0y0��$�fIj��RD�mK��X�e|�Rv,�c=�̸��g�n8}l"a��QT]���!��{��;�Z6��7�qp�ġ-vU���84��+�ͮp�Z*��c\R�3��������n��q-�����Vc�]֣X��ƒNhE�x~�E��<lK��pe��%>+���>+랍J���'�d�dhI�9l����j�Sr��J�{|�;s�R�����	pa�����r���eؐ�N�w.v�UNi)_~�Ll�ꬕ��m}��ɲ�4���������j�4��?M�����:�G��Ho�i���) ���z�ᵀM�`ң�:��~�ף(� Je�Nm�v��
oo�{��|�,Ŭ�I��4�����X�޵JtM�Q�m �/�)	�8�N$W�#>_	/�uu��.�ޭ�~�0���h�E�N�q|;"/�X-J��L��!��)�AG��ڝ�)��$���Q�-[[o'>*& �,U86D��q�&����b��	�M�79çK'3���Ь8�������������Ƣ:r�R�Nn����!I�H����X���gr�0�$�&f�ıK�0+�(G�oS�C���Kh!����9ܯtʥ0:ۣr��ֈ���h�#�D{�lъ��6;���9}X�3��KYO[�9�Hb��]gw=.-��.�x��t�|��X�T��b;)'���D�{�C����5���_��AR�Aۺc_pER��N72v�!r�!<��1"��2a�_��3?�pX�j��B��GZ��K��ֲ%�Mul����2�_����"ߣ�r�b���H��6LkT��I䞞8 /T���ʘ��Tx%��X~eʲ2��<\��ե<��;<�\���\"_ފ�-��G屝b�����GVU~�c�`~L?;n�Ӧ��7��
��k/J� WL���7w)X��0D2=G������;q_?����5�>�_�����p�xV�a��Q�P��8W= c8܎�Ŏ�X7�I��~�ko��=�nr��ω�֡c8�׿�2�k��4�B��@��@��Ȥ[E]�-�gO�L&OGʁ�[�L�qՅ�
B�m���^�vB��y���Vi,��"�2k�$H���h��m��N[�0�g�m]Z�w��!���@��t�6[��v��ᷝY�)?s����[�'N�3	��s���n�O-�$Կ q7+�o�/	{m�P��i�yxo���Z��.1�;�<B��� wv��nT��_�h���jz��B�/�]n����G���71L���������/�ޝ��"�.9Q�suM,O�{$.�0��S�oȅ�ݪB��6Z���]&FH�y�D�j��n�_k�`��Qጸ���T%a��	Q���3F�׼��*>�����m�sR�(�yA,\��#��;[�v��&�,��ig ���SAx���'�6�q)���ZW�ud�F�������3"�QB�W���~�m�{1�=���=7k�,���<[����l>Efg'�"���3uR� oݛ|ꬨ/8l�-��@�^3]�nS0a��~��C�ҵӏ��,�LH�9�X���X�ƙ��犗�W/5I�����+�*��<N���)70c6 鸓Z����J�H��v*��.��Ꚗ��Ac�/D��@oF�md,-W8�����c=hL_�#�}�R�z.L�"�ќ6��5��w��W?�e���A�.�H_�n=s���V�L:�Zn��r��+u�Ju�~L�zg�i4�ג����Y~�Ŵ���9I>�z�<p8 �t�k��S��u�se��n��r��?��	USA?�(�i�%4!|�v����^�E��%i�k:l�gHsu9H(V�Չ�tDp�/iF<T��>�BEѷ)Z0R�[$9��^p*Q|��ҩ��鑖J��<wirD4��^��pk��t��k�G&�Ͽ<o��:����T��=���g�0�$���i[j��P�z��porP��	R�b��/�N�4�x�}٩\a��&e,}��"xEvpQ��I���9|���g}u���sOWvI�h�M�/r�!`�f��`��m��P} hC�5���p)*�����i�k�5WwH<�`~�)��qi�#L\my*�໓�?�N����̖�c���ɳ{A��1o���,�WU�W��b�e:��-�������|W(��>t�~���Q41�,��%�4#�V)e���y��J�wٽ `16�/r8�@ŵ��^^��v��聘fQ]��<��#w�.3p�F/��z%CKZ �� �7��_�#�&��ʉ��z�s����q8��e �^?u�l�7)TX]/�*�K�66|m�91̓� ��������\�W3$�a\��VI��p��=��9f�[�g[��"a��TX�s�,[�Ʊ���̃�C�嵼��K���{{-Z���J`u��
�#`�o���	?V� �C��\�/�+��H�#�Dצ���*�zwp�z�*�|y�;\�E������
��˸ܧ�o6��H1�b��U1}L=�$8n�����99����*'��W0��+8� ����b��jji�jY:�1>r��>wr�z�/Z���0Eo�t��?���,\���`m�"x���K� �*�
�bK�$�Z�Y;��&Y716.������$�٨�n�v���	������81�Ĵ>���-��*Ӊ3�$8���ܴ��z�*2��DstS�:3?|zvʉh�`�j.���Rg�t�!�(2#F�z'D4�"���ܳ@`���yƝ5���o�R����{)�)$����O�ٲ�k��E�\�<d?�G����f���u�m��Ӏi�Tz�U����'�1y�TB��Nێ2s��GklN�t����_%�.���O�;4��*���Rf�;&kf�|Ƿ��T^��f\~{�����ryx��s���*���ޘx"Akyw�O��A����u� ��C ���r�ʢ���(r�'��ՌY�A�)�Y|QEb��w�������U믹�ʏzU4���6�o�,�6DVk�Ni) �	iBv��/��nO��!_>�5��P�HD+o6H����@������� Uo��+PC��$����9�����xK�!6��`�T��E0?1pd�;����.�/�[[��ɏ���i�xv �c�H�qZ`���1��+��� g���mQ���6~�*{˫o
�	am�OYX����1U]�`���OZ����Ф�Vh�e�T��@�x��-�4X.��Lc��/�������*V��x�׶"�k:��Y������}"c�ˈm�C�5Ǔ4� \/�6���W��Aj`5��? �,�+ra�T����2T����*�cEz�iOto������G�!>9��%8��M4���FW�~^���>Y����Y��,��M����!�����*2��x���Ӊ�$}�`���@��w0�\�ăg�~5�{�J��T��)���.D�,G?-�����_z=�T���Jo��i�]s�r�94���a���B�v������BmF���' q�]h] \m��: `]����K!C.���F�F>l��Ǜ�H�P`?��⻺İ�{�+����ߵ爷�6lc��Q�լ�H���ԍ>v���`��w�~}������,����~����L��,R9z���OG6o��"n�@(7��.��$N�րW^��-��`�'v�:|.l�4��~�x��H�����D��Ȍ�Z��Og�A��`�����jas��%��L��Q�EOb�W�뷦L�1���'�YgJv|�$�?�h�.K��  �Ϫ-p�jy�80�^7�K�|��<��]�Wֳ|�H��!Ŝf���L���䷀f�a���\X�֖4��/H�i	Vs��f< \�m ��x)�Ǖꥤ��g�F�y�o�0�v�a��is���.�`|)T�B�E����FdN�V�۵V����T2���y����a^b��K�%+��S��Қ<_0c����پ��H�@��� �8P��B'45u�{3�h��ms�4���\C ���!�e5��U.���_������9s�ܲ2�X9T�S�|J�P3���p���/��_(��+y�(������p$�y�?�߿�X�^ޝ,���J�ձ�V?��_O�ɫ�F�;s�>� ��� �G�+��U�a�5�������	3r��N/em�Y�B����<c`�!�3��F�"�r<��9�AA�����~��z�M�#-H�-���q �F��##��ޛ=�,�2+�`E(fV��rWJ�G/�������lU��_�(W5_G��_�q����4�����+S��i���ey�ϓ��C��ڃ"��(��$���-e����z��B����	�"��!��A��V���L�ʴ���:c*B�0FD� A�
���X4��s�[&�'�	P�J��d���{-�W����	h"�A65�<�>\U�z��~Rl��6Oe:*�4Q�#����O�����)@��bŠ��M�^s���39��^��ź0 w���籟7���U�֙M��Φ��?+�v ?�7�Q߽1����u$�I���1+��$(�F�T<�L�9��7~�^~�:)*_Ҙ�?�Jqx #h�萮W�]�Ԟ]��z���6��DCa�nS��a�r�|�f�Џ�e����'e��SͻT�����Ο���H�:�7a3��)XT�B�]�%0G�Nq�̛IS� "�&_�UZ��EΞ����p6����O��#�����Ν��=�Y��9U.�i
���l��FU)a%�8����S����T��6z uY�)m}	�9j��1 ���$ìq�5�?�ϹUˏ�k��M�_��g��a�[�����	e��wz0�'��ɟ'Md��۟�^�ԥ�=/)(��Q���w��G)\4D����P�����_��� �y�he�V�9o�Ħ�ɮL�O�Z�a%�?%�j*��gM���Tsy�@!,��W�a�T=]4]�����+�9qW[]��$k݀�}��.�g���ײ6�������Dz�3۝:������a}�exV�\��0��]��'���}!���{������-.��5�PW[ː�QL�/�&���)�H���?��p��D��] `����&�g�+���w��n5�/´k{�r��p�Q�7�3�~�� z��P��Q5̫8oC{�R��!�Q{"�V�U�޾��B_�qǫK��A����Q�Znӵύ�P�d���=�jP��F,��AN�nmh�j�C���톸+c7�ƴ��t���������'�lH�[q��}��Rc.u{�� Dk�7X�<!��8|P�0Qz��Gg��%���E!J��iAP6B�o*�����i�B幹�TK�Ry�^�nQ3i��6��B�X��Ty����P\��|�Mō�AFi��I��"�󡑋��ܞ�d��}bΟ��X���20Ɇ0"<��3�p���m  o�����Ұl���$s�����>����iq�O�I�Jg2�3*������K���@q�"��Q�$�S�ſ����n�9�O>q�Z	�a�?�s�M�9)�O�@��	�q���B��]-wT��c�_G��V�1�{Pa*uk�#�Ee���R����"�����u�4�[�[�X	�c�q����������qYk ��o�������4����8b�ke���#J�j���O����5FRlJ��ԑ��th���yEer������٘��x6~�n���P�ۣ��Vs��՞"4�%�jK �Uӵ�����?�k���+�n�����R��Y0��*Gr@߁�M���j�'U!?�d��4/?n&�|�fm�@�Ɖ�
T����L9� ހP��	%����ESw
�o8��$��a�Gqb?/�{�,TMU�s/:�[��[���	sM����~j�g�Gt�1{��u�/g��1o�-���g�Q�1���4}��G9rl�Y.
�0�I��<b�8��〹�pf��HU���ʢ�Q�I��ܦ����Dݟ|I�,T�(���Z6|�A���-/ޢ
,�{���1G�  F�}�&V,*A�F�S�b�?���|^�����oAݕh�(ABk`IC�,'v�Z��0a�N,�v�*�E���z^{�cg�؋�n�͠wD]�@�6W53�A���N�8���C��;��ˢ�W���v���!���7�n��(w軅V9Av��b�T��|���D�������Kb�zeb��G|1֒���W�Ε��(ҷ���>�_/m s�u��8sD�cc�0'�ʥ��0G�z�W�ʑ$���&�	�	O�x���}��O���M7y� �S��Z��s���wiL)#�S���6l=����>Sݼ<URc�O�u�;_de�"B�"�_y���6H�y޾WQ�n3�#N�r^����rT�͵q@럗A�y��)��b��rXDF�1� �BmE���������Z�� ��ty�W���&���������>3#�XXf�JIb���j��nu;�W���
��-q0��x��'��wdp�I����*�O5�8T���4���r�J?���q�$t�ŉ.h�t�
�.��G}Ǧ�ز�9+wT8;�h��A0���!K�B�׮wd-9���]ݣ�X���7�
 ��n"��R8�<O��tx���@z���#4��W7���ۯ�΋u*�<j_=Z'�iiY��:B�vgm��4�#�%�s��t��y�a��[ҭs�dɮ�P��\��� �87̓���;#�c9PE}�u/ G�2���m{�s_���Y��q9Cɥ�iKVi��������v ��Z�wPԤx�V�{;P_9uGL�]l�$Ӈ�ٙh1�ц>A�rR�����X�3���4 �����D�i���s��Y5sX�<y��O�4 �� ��N,�i#@��`p�|�n�$�<�e��%���3N�ҷtShw�v���>P�(^��X��H|�p���r��s�`	�N�
�t&J�g�NTң�R�)�\.u���д<��屺��]���cl�<�U5�g^���YM}��4zV�"���\|�x����t2_F��J.����
�Cz:%	�<���;/ɧ�����\�Z�����\�fk`����h_���jyo�c��#�z`=��n�÷�"�$v�p)�P�vA�tU#Yu���*�C�������SG/k����~���cfJgJ���2�-�Mɞo���n�o ���m�dé���k�ſ�$�yucƯS���D0)D���P`�{d}g�3�z�Af�+k�SfJ��~�&G�ڽ�%�Y �W��������5���f$h.h��4�j�f8Z�U��糷q^m�/��^�/����U���J��Cڗ�{�K��<��(<N<�A��J���Jh�]���/��mk�5CtR!�D;k��b!��3Kl���s���Ϗ���c1��b\���n\ �S����K	]0PF8|��z�r�F��>�m��RA2�R�(L��e@hVSۃC]G�����ʘX��%�.���'��������n��.��Ãw�r����YS��=�h��y�&ɕ
��PK|>u�b����kD��%�^�M��I�������2&��"n{��E�4�����s����7��-�(X���c���VxG1��_J:V�D�����o���;��Z �X?���W��~�n�zi�}]�>t��_4�e�� �h�˪]�z�����ے$��w��F[*�@������R�*��$���CUh��!��`�=N֑0_- �ci&H�ƥ
��"/^l�9������@��T�3L���_s�p����g)
R^�� 
)י��3l���]��v*qS�T�^fb��;��3V�7^r�����u �&��Ƥ��V�&o�:��Z�O�5�ׁ�8�� ~�+�����3����������S����6Ժ ���s�% �;8m�[����.�4��	�;
n��o#R
����s!?���V�����+ľ��hy����#�^�id��S�w��JLJP�-�{��L�v����f����F��E:������8i{?�`eL�мZ��������<�A���h_�QR�� �PB��V�)�v��7�/��d-�*��y蔻���⃇�B˞HGCN��ˌ���o��R�G�d��a�'���=GgCƊ�'��*�=*�p7Vc_)�4b�"_T�� �1��PR@�����#	�ou�ָl��0�.���rf���B�Aͬ�Ȱ%��9y}��J����UV�ZG�S��dя5��i���a�·�]\�'�����Y)�Lg*L�U�T~�	�S�쒊ǌ�E˟D<�H_����xf:����3/�Ř��>G��kh���F���y�M�n@d��Oj^�·2�-4�>�F����������r��_jn��V$J;�E��"/*L�㺻��s�^���q\Ϭh�
b�yM�CL�M3�e���mg��&g���10.��9�h�q@U	�?:�8)8��)Wڞ=u����kX��\}�������G.i���[4�c�?�mҰ�i�\��R�������AN�v_$�z剟^�(s�8�W�,Eq-���.�H��h�u����� �T�m,g�=F�{�#���p�<,]�.�1{Z����U�:�[?w㱈J��X�f�a�U���͏��v��G�\ל\!^��TԵ`��g$��@8[:��Ǉ�
��?�I���t�͇;_�&ڲV�?>�����/�ㅍ��O�D��.�7}�p�����a�A������(tNP��|U�����#��M?bJ���?]�����$dNFaz���i�%�����5JG����$Ndl���*�x��0�{d��y&����@���娚�ͩFJn�,Ze6߹x��n¿��m�\I�B��)��o|8�-��~��{�&a�%�#��F<���_�Ҽ���Z��]~��6��}<�}�}b=�x�i��p��I|����MW��ѣ����Qox���b=z,x C	U�z'Z�={c&�p�d!~�p�X{v��ތ{NZE�;ڽʄһ���7j��7�"���&����͉bt��!x����+���$�pM���, D�I�&�KK�#�~��w��7Q��͙%�˶r��f!}�����qE�<�F��Ԟ�|�} ��-M�W�Y���cFZx��^��|,�j�y���4L��`P��Ƽ�F�
����Q�ԑcܘf�W�r�|��\�����#?H���q2�9�e)������ⱴ�o%f��|�0�8���7�䗆�9=�8���y�z���!�i�oF�G�Q��@�m:�1{��N95�)����
*ƹ�o'���uPn.����N�����e��$�︘{�;���|�Nc�#��E��� ut�u�|>�he��Y�"���p���\�B�:L���F�xe�s�g�����i0Z����\��"-���,1	�J���]�/�5>p���B����b����d��'��IuxLg�X7���ʴ�
��6�Ua�`�흷�==�G:�p�6@v�ƍ��
����8n<�d�Z��"B�.���;:�(�߫�����bH��1+���MD����W��c����f�?�G��-׉w���X_\0���g�Q ȷ�{A����pM߹F�:�^����b����(��R�`B�O �Z�`����$C�xl޼��v��׎41���+��|�o)��'1��T���(RXX8}/���n"��^L��1�j�!�j�����Yl՜ƱȮ*u7{��
zUC(2����c��g1xF��	Έk�s��T����2��З�_�=�m�S`�K�c�ڍ]�3�M�#�͠]�n���k��,�R�Ǵ��R��́�����k�Q0��6����U7-U�� V[�iM�v�����Aa��e ~Jژ����dd�,A��m�"�����x9��#�׎|��$C�uٱҠ�Y�yS3����F~~�r�1��|Gn2���T޽�qlk�Q�^��G!L��Bo�;<���ql����0@`����t.[��K�9���&7���iz��n߭�>1'�/�0�����!��Gx�8�����<����_��Y��عwB����)W!����J��m�̼�@ٓ�V�w�����$3u���ԇ�߿�6T��QL��>��_1 ����GX0<�
��@���-���g����oZO�D�ߺTJ�M�đg�:��`9 �spz>������-�o&u�]��;8���6�ܨ,�?6�8�m����{��#�Y�{tМ�82?_i�p�蟯���
����ٞ���˗���:E��y:�0����?X���\�[PXm��ܰ5~��}��;}��~%+$�p��~@�22���~7ba����Fh��a��2��H4���9Rj�WRu`y�8Ŝ9�5���cB|3v����[`Wm�u��������q�Ƀxץh�K�v8V�Su{Snp�p6E����[�qw��p�
�l�_zy� ���^����k�Xx�R}�0������ӕ��=�#�f/�A�>�OU"��y���p>p�G*��� 0�P��y���9��4#����9��������E��8���W�/+wr��`���C�8�M�O���'=2�Đ�H?� �qrf�F�}�-`S`�uh!�`O�-w�#w�$s�
ؐ]�a���6L����K����^�&i�ۉ�16H2U>�F��
�!�[G�^�M�;�ÚC��n������C��@�B*%��!Jh�ob��pM�����}��V��}�\� p\F1����M��K���'���S��h�J���ۭƱF������{���N=�8�zA���թ�+ao
2�^�3cG��g��/-v�n�`������Jü$v�T}܊H���$g��;�j:�Z�Jvaz���lp����)*�>I˸|qmoLV2��3�Is����q�rc���c�.��':[E��{Oɕ��?p�O�-%�f�/�b�J��B���tuis��<��a��C�~`~�ߺ¾���߸�} 04}�m�v�_I�c�J���SC���Ō7m}`��P�$��Q�Q�'J�`u`ãI|�_���U��ߩ�0ҩ��:[�e�AuVHP�w�z�殅�U��E����=^}�G�q{5χ���:O���ɤ�?҈|L�/���5C�z��Sh������E��/:l(y�@?_�A1���A3\sU٭d��������A^�G���Dݭ�h�3R�������!�%���+������� �mKo<��n��x��m�0it\"ׁ�<'7)����������,����%�5�Hg�D8b�'���a���˚��_E�'-�N
���/� ���f�nH�BNUk����&������������8���^s�Ce��9ͮ0.��a�j�K�?;ҙ�QlʳN7�
��-��(�7KQy��y�2<�����
J��_r����Xo����$Ua��/�:�_9�7����D��Ϭ�y# ���L_
�!��LM�R��GR��Ȥ	��%��?$��QkI+$Y ?F����s���ۭ���[z��L��������pJ���������8$<���ߏ��@���zȏ���/1~(��9�8��h�k�ƽ��bE���dk�e`VNQ�^�^�@�S�n���
>��V�?��2䉴����Q���p�[���ف�-���̢RšMw���;3�(C� �%��u�����j�s-�t�����<�PMJ�K���ep����bVA�A,��ŜV6�0�u�@@e�3���	�ޜ�9��Ξm+���A����59�ފ�	�?��:�����N�[D��H�����"2�C��0A�#E���!!��$ҹ�=��}~{<��ι�u]��>� ��(ĵ1���	i	��}���Eᇣ� 
;��֡'w��sc�/�)��@(�Vb������\�����lx�1]�\9�ϒ``���Gޏ>S��v[7�"킰�i)b�d� 
���z��J��p]�|U�~P����p��k�A��u��:�ӻ"�D71�����WZ�N��Dpy�u+ �a�#/]��p���6���ܱ�Ze7ױ��M�����90؋�ј�J!���0=��Qʒ�b��K77����e�9�����[���� � �_� �~�q���	��f����b2.6�_/c��s����钺��Г�9'��<�����${? �|?<*����"q�+���k�Ҡ��L6~zy^P>T���".y�U��ч����ӻ�:���^�F3�u�i	����s � 	�2�`p��L��n+;D��|@[=7�oеY�KB+�1�TyM�I�T?���cE���f +�'��r6�qw�4n��ު�CΛ�{h�;2���3Ƃ����x�af�]�l�F��x�O�n�a6��;]���^VQ�;c��������X��*=�l����P����Z�.T�'4����o��.�}��b�)�r��l�%gk�V����?��,�K�l�ܓט�}�z��4A��g���~轩b+��z��
?��P�^�)Lt��w|�v-�z�?�Z���[������>9��� q��5�ԘǑY2|�At�|쪹�Г:��U'�8��)�����3ܪ��S����ò�w���E�|x6��l�H����4�[źڹk�|�u����z�����$Q�!�W�|nn� �&�-e��눜6㾡��q�������1����K�}7������X���,{~hY�UR0�hrr�i���9�j�GA<�gqӍ>�E��nǋǘh��F���K['H��ro�g���Y��G[��󥼢�ϟ�~kq)�hadd������!��m��z�ES�$���/��.�����8#�K���qi�;�y+>��O��2�}�c���JfŬ��+�Y��!�f���C����_���Y�U7�@�T�D<Z���̉������6B������ê(Iy����2��?�D~�p��z��F[����A���i��Ɓ��_d�����X���Ŕ��JP����km���D(���B�K�	�+ͲI$��[�_�\܍���h�
�_K�2�ttt��BiU�d��7tS��yyy�u)h��:�>�?����A2���m�&�a�S�xoB�9O5S6�j�����~����є�!g�_)�������p�x�0���6�*:��%�����~�~�\���:���븥�&����e�a�.�ߕ]#�4�y����ՓH��"i�d�)����5X�6a/�`��e��ÿ����>��zvq�#���e�1�X�f�k�F�,��\�e����bx�Wo}�Q,N(HF"������[K�JA��h������z����|��!3�km���_����p����xb�R����0�~�b��a]�ޒ�
�=���'��g<L��/"��+_�/���.�Q�	:���Q��_�S��Q!����cU3�����*Gf��4���U��?R�bw�FFF��}w��$H:Ii
��7�#ͺ�jB�<K�b�j?;�_�#�?^+B�D��i���}�B�k-B$��_�iR.I�(�{�ҿմ���V�"{6��l��hb
st��wQϚN�
�J�ĺFAUT���1��o[�AUb��F��c��̸'�J�ד������Y:����DxpW1	ZS6�%������{s�ԂA�����?�*0E�Z�`q���)rj���ng�O�ǵ��[��{l�+����'�����z�+���<����|���f���~Ǘ��xI��VS��~��W7˭����w_s��V��]B�/5�P��QH��e*N�e)���	䢐���n�$����I�����\W�!���%�ө�W�3���w9��[�d(���;G�`���0�g���1`<��>���7$����͈9~����=���L�����R���M��A�N�Z�����N�H�a�u�	��C���h��,��n�S%N�rTIߋڄX�zm3���wj��̼��9����7p����x�FȻ�XWa��xhx�`��c�R� W������j�yc��DB�Y��mӭ��9�w�2�VU�9��F�CG;B���Q��P\]�+���=|L=�}t[@b7���L�����Np�g��/y�5iY)9�����;��Mq0ز�9C���Xp��,.���*	t�&3-S]�Cun��*.�]��̆F�>O4�=w�r9ܰۉ�T���T1��,��Ӕ���i����%.��`��Nʦ����ż�ՎG�ܪ�ݰg����pҿ�mA���@�'� x�=��}5�0�/<U��O�2�jJy�������|������M�B������w������'�o����(2c�G�ۯg��w���솢s�@i='D�B
�n���o8�U��%o���w�~(� ׷Q���oź�v	�?Z�Z��������b�����K� U�_����{�˵����zuy�΃Ly�V�ۧ�waRV@a���4
��T�QBp�Ŷ���(%ݡ��I>���@>��P�y��^����뇡��s��_��w�%)ͯ�$Q~l J���-�چ��I� b�f�byW�s�r/�/�����g��C�|k��v�V��e�K�F_e\��%xz�G)|S����ĸ���[���tҙ�ǿX��~���2��;bgX�L�9�yo�ë����^0��ݪ��Ʊ� ��([n��F2f&A����o��BQ,���U�06n���.�ьxJzٷ뭉���C�q����ǁ�D�⿳�;�`HS#��	�b��qԎV��������xO�,��L�������iW�k��Tݜ#ʕ�z��c�w�'q���tPN;y�T ���ϟR�%0X��W
u��\`�G��U���=�L-i�l�/�M�s�x�4qH�&�{��;��ҹ������0��Q&9��r���3�����i�G�7��V.�	��g���~?��:I��q�=m2uT
�u���1Ȝf��N��M��L�|Զ��-w	ձ��������m�_����W��+�,�'�%i�ư��Y�G����]��I3-��JKj��}Pxj���Uݡ���� E���a#���MA�*��O�5!W���0��I���YI��^g��q�2��"�����)�D�v�\8Q�7��%U�#zU���U�|�>X:�3]�'b�9܃�Ҝ�x���3W�,�����fҀ�տ 0���Ma��Bls�~�.;Q%����ď����zL#��C���;@|	W����i�j�`J�1e�-�ϓ�!��%W�o�Af'�[�P@6��K� UYU�c��dM�$)����H�.:,��߲�G؀`6̼���i���dF�\�^�YQK�B)�>��F����T�����~�.1V����kޣoj����',��،�=J�Z4W2W����	(X跳�������o���d���f1g�BV�:",�E=>e��rFv@�rڀ?l�yh���5������P,���%0��[ȓ��텴E8�Ͼ�[�/&0�F�~.��A�u2�]�p��.�4�;��cRH���Aa8��q�ke�:�NLV�K;(�RW`�ՄDG1��G7e�4&/ED_U��<�%��VR�q)��|������UɅ����
|轠�M�� �+���{$ï� �-��ڒ������/�=t��xA��V�̽ioO��\gE��?�GV3%d���N��Gk�/�ӄ�Fu���m��劶c^�`��k� �R�|�6���;��Vb"/��;A����AX,�K��_��TP�U�?�ܿ��<㪺�L�/�&�k�T���K���*��;xQ�`��5{�9�-�������9ݿW�v��X�ѣ&�>Z��+j⡅]/K^�%�\��Q��#0�
�a����(���������إ˴\������  ������P�������e�����Ʋ�0���_ϕ����/�Id�:��*���ٽ.����Jn�?�|�i!D0�$pk�jn34���H�
�?��}�Ts���AS"�I�>M�D����W�4e�)���Tw��[�Ά����&@<��/ؑ��kǿ_L�v���Z�"q���s�椛|MꜢ,Ro2��b/�\2hy)W .��LB\݊�&R��3�Y�ן�Y�Y�a�9�F9����_����M��S�5��9�M�T�f�@Q���uҵ?�(2�p�D��~_�
a��Y�Ǘ���� ��������(2$ȿ�5��=-?�$� k)�)G±���������+��X1�c�ݧ�,�8d��ȅ�fn��_ۙ�1@�C�cdܚ9cύ@����)�2B�2�zB>���):7��]�a��L^�))1��;���2s�tВ�͛;��]
/�2��n-г ��� t��P ��J��+{��c�5��S4��1A�U��+��_�I;���V�tɪr�*�+�aU�w��\)ubSS�t�	_ی<;���<�[�H��4�&(5<����8�j����H����� �9q�Ϋ�j��3/�L'�E	I"��>y�$�]��_�,*i��J�)ą�K�q�um҄�I�@�oN���\`E���_�m�VHEN�V��T�Y#5c�~�3/�΢��*hg��ފ�Ȑ�#5WiMaO�e�b�4��te��L2P���7�����@��D��3MA{\?��s�)%��c?�\�C�y��}�'��#S�����i�)���?{#�>P�
#T섀}�~���"�-�}?����%�?���n*�dw�v�wb@���"%��y	�P����^���r~�w.�f�h*g�n)+������x=��:c���`�_�����7����q��7��k�B{���?>�)c�9^�m����[��n��d���X3�h�ә���� u]�ʙD'I�B���%S�xī��K�;h�'B�3R�Aن���P�i�~ _��"��t���'�L�
f��ontڏ���:)� AzHn�5-lD���)���j�g������2(y���y [�� <$󪜩�.쎳O����a�5�`�m��APGe`m�R�R��|�=8`6h>�Je��.c �P�[4dI��" ��\"�xݍ�|�R�'���<�� ��.7Gp�ܲ~q��4#��, Wվ(a��*GM���_
TXd����8�V�i�}K���<*n�S�T�0R�"���S���Í�����T#m��P?`W^B�+S�������o��+����L$����rN����+'��<x�\�D䢺�O���?���6�V�O㘸˻��[�;a��b(��h�ͻ�C�Y4u���[
�R�}�z<��*^�Է4_)4�~�W�g7 -E��/:�s�"�b:Յ��J�9�}��XZ�5�aQr10�������/�fR2F���v��k��L��U�M�*����K��3����5����k�"�5��܅�/���v��u��)�w`Q�(F��a��M���I[��<?�l��T�����GG�k���n��������t�f)�#���y��Ʈ���`�r���f�Q�`���Y�3Pb�w=Ak�@e�~�� ��)�̑������LJ��h����iT�ӏ(~<K*�bU��������	Ez����;�g,1�_�4�Z�4�6+�QQR��*?`��d�.�>o�fC�7����_m}٫���/)��c��q��c�1Pmy�g���Q�U�IȲ����Ε~��ƞ�QX!���2ƕ����]�i�*(wl�a+d�؉�1�EN��[�>#K��H:CB3�"P$7:d|��y*�:�0��V"O�{㝲�-��T��7�L�;,���LQ�f��K�Q�'�P��|��g��t�@b-�{�3�40�fwg���Eҫ|��-2�����g��m�;��{�%�8�BP�mR�D�cQ���y.�o�c�� �\헿�`�ׯkl��
L�s���g��V�1wv������;ʀM:QO	��w�������HN1��c��F����Ay<T�����6�/�*6`%��M�+|'tu�,Y�H�*��Uugh����'��ӟRS��Y�=��}x�|Ô��G?�=�w_���nυD�(���7��o��������I�m���2$�)w�Z���=����h����&�3EO5>��4�!������|k'��_f���$7�<����f�	:-���Ĺ����f~a�ʮ�s%������ �mucFI��ɑ#M�ծ�v�/z~vo'�⥶Ĩض�zK`.�W�)8���"�*���^}��V�@$�_��?���d[A�Ĭ�%�-��}��ψ#x�<��~?�y��� 'sn0��&�?ו�`_"��Se��+f��ة	�yʷV	ϮG.�Ck��-�Q�r��i���[��e����|����ٞkw�"�g��Eܿ��*2�8JO%��>���Сt4u�������5`w(�z�W�[�t�5c��8]��XE�-���:I��(y��mv������r]��X�3�0l��u�A�(ٿ@1ya���Q�F�n�Y�Ih@����6悒kEd7��s���-JK ���ш78���%���VPC���,�Q5�?�LXq ��"�A�K&���]ؐ�U�Ʒ:�&,�n7	o�y�,1Vx�dt�MJ�KN�ʏ$bI%I�H�+��=łA���L{P��.�X�������?����gI�L[�Aos���5Ŭ[����_�zY�W�(3��y��w�R�k�ːLZ �n1�_�M��Y�(,��Jҡ��X�Z�woX �hBQ��jP*�}�7�3i;��0YI��N��ɡ�|(Y�����U��/��G˦��&Vac_>AaU�l���W�5��m ������qhs���zͨM���Y���l�돏ꚾ�6�\=���-�y_�;{[@�:'������8 l��e��<0������HEN$�Z��.H+�ʜI�H���`N�S���/b��H�&�	�蓯��<d7G�#T���V�c�d@c=L���ί�}�Pϓ��-��1���Ɠ�� ����m�SQ�a�n�\w���"T�@�O�Ea�\"��g@�S?�Y���1�:O#i�{.�������FOq�&�M��Y�^Y�P���?��?��������58��I*Ky3t���|��Y$�Tja�>��эo�NO��a(؎���뫎��h���gB0�Z"uQA ���aY��ˣ�
�1�B��d�:�.���nRٛL�������z15Qv��2N�Ӕ���������ߒ2G�͢0��
�e��2�c�,�l]���g��Yc��^���c�L��:�< G�N"���e����g/���(�V<0P�6�ȭ	! �* �:B?�/�Yv�X��Ȯ��� ���J�c7������T�)t�f�u�h/.ٹ�6���,��$�ق�@a��Z��ŀ1���N��M�x�:|�Q����6r�e�$#�j���W3/P,���S��d�j\����|�'�eݔn$��Z��N9\���\`/��]����~(���:�4�qp�zx�x����1��F�,z�EDF�Ւ�Y�"�
�h�>�d2Ql�s��=F��%��}���㠩�_��*;�VE�rGL�/��#�K�
B��`w y�4\��D䈩]�%�Rfa-}@�͢��,�3u�,�3̆�s7��ȕh����&��45&�)2�n!xa��=51 �td�+�T1�ܢ�~5ˮOp�0�حO<�O<#�/&uuf���w�҃G05���iF'~�hV�A��%K�:_�ۈF�ݏ8��ȑ��FJ�A�F��� %'��6&j0�{���51�ȉ��B�x��Ci,\�y�a֋��
�_��Lɺ �?�V�ꏯ>�P2P��oW�ŷJL�O�q��h�����	�P�I��Y1裤ܰ�(��von��������5UK��~��X�Ăa����@�nw`�-
,<j�wC(<4��3p�L�� �~�6.۹��`���������������SZ�g�)�|=,[��Bj����!m�36y��KS�4��V��/��.��)*{2�����<?�MQBW�
��t��=��
u��S���Yg���HM� '��� }v`����8mc�He?{����1���įt\�/���F�C|W���3�G%��6ޤ9�E�k��_߾���[�p�o�k���O�N�&��P�+�B	�.S?�a�P�P�۸>�{2���x��ck���@�f~��H}��٫�	�u`߼�-^�q�9y@�<�W@I�8�N8ȴ"雯�>9�t�/�nn�g����+��1���J�ڀ�]U��0H`�����C�SRp��.�����-���-y�+q)Y|�D$��J  r�s���E�<��}촣0MGK��oTB�*�oW9<���6N����6�F  u�HdT��O�6�ⶓ�֍�.�����G�rZ�=2�'D�i��e�E:O_���E���Iw8F~1�(CD^��͠5�<M���l
��`I�G2�Ѫ6y4oR-�G3���{�1��c_�P��z�/�:`lk�!Mo��i5x���1����E7.ŕY���d�T���v*~��G��y�`rW=���*�Sj4;/o9�Է�\�[���hB^q�ح.���F�J^�?)�RT�L�(A]����!����)T�)<)��T���yA��k�|Ծ܄������4�m�����@Йox�N�c>Ŕ/�~O<��}�3�T0p�M��۫O�<����@�шՋ����Ќ@��j����·:q^	|��0�����	%�y��D$�=a]p�]�*틵 d�A�9�ښY�1��|��K��}L;'%�Yk�'!=�F��̱��C嵤A��y;t�"�a�E�Nzrj��s>�
�x��c�:<�;��ɣ�\f��س�HA~h~�8����OP�|vAr��i�&{t"9�q5�g�H�|��A.��7�I9��0Ttt��f��2�٪�����7�i�L4�Y%ًyB�_@?,�`Å�&�N4d�P��!�1���6�ǔ���ksl���7�lIЄ�!Ӯ���n��U�
�*8�A����L���s��D�Xf��0����-2���R�(�ᖆ�~�7/���X2Kj w�6�ct���7�c67�8؇��Y+�����4ze��0M�����h�J��:�	j�P�oyף�d�|�ܐ?�s�s��~8��@�l�W�����K��g�9� D_���E�l{@�C�P��&��n(�����]P�V:lj�J<?G���ˊ)�����;W�W8<��LR� �)��7/�~<2�4#0�[mx`%���G�����f��v$��B"#c�;��M�}��`93�A��A�@�S��ߓK�&ޑ��e���qO�˳<B::����֦�Izp\��W9���v96��k��;�{���)6נ��'�+����s�"�dj��oFe��o��>�v�[ی�Q�����Q�J�-��}?Q,Ƹ���k�5�z|h�#OV��\	 y}P���r����ś(\�>�\�8�E����@.W�w����e����yمCf5��ܼ���L�>,�~�� n�\�É)�MF\�YQg��R����;.h��(�[�~Y��/0?}
T.�M�c�[��äs$�<�{��0�e�����ZU8�/$��1�>��];��s�6�l��X�X��<͌0�)���\	ǰA?�xD<'T��Z�U�&ԁr��Ϯ聫:����,�����p�b��Z�������˚eV��!�Y^��f�=[ E�h�<J�]�����-I�����Ѩ�	�.w3x�-�o��z�����`}��@)%`v���`�a9�o��f�c�O��i!���7�3t��UD�xk����;mf�9(��e�ŏ�{ט0z�";޺��@�3N{G�}�1 �F&�ix#��j�� �B	��D�GnM�#�p(����y�K$���C�LKy�xp���(!2{��[>��c&�go��e�j�$$Hʑ�i�z\�4pU��C�B����h��1PT)b�"���yjO�n�,S��*�y��Bc1�u��=�)'��֍���O�����m(z�}<DB����X���т곷�kek�}�=�0\�Z�M����+�MkUp�G)���[�w�H��
����eU9{�s�J �Kk=V�����T@���}Z:�
/�t�6
��2������V��h:�2�������I�S�����e`)�q؂	胠X.| �6%�[z#s��HG%'3l�a#�"��%t��l���Ѱ���`6MޏW��g��窞�.�^��r��|�L$r��1�s��_��@A����֜��@'�+· Y�M�%�w�����2^��c�{�"A��m���봓�����Z�Ax������L�q�������Q���*�-��%3���A;cqU�\�A��,����0Ѷ�y �ʕm��!��:�Н�g���u�38����W$�_�G�U��J,��@��2$����g�&�?�����d�X�UH���iHuF��삒�U�ʖK��˫�_���-����B�/v!>����&2r��� �+`���.�,��Fq�N<�)R2F3� U�Yo̵|n�r�#Q��CU̴�{��ݙi�j�_^�C�.�ʒt�iacj��̀���O���l���e=5�� �j�����<���<�)�j'O��1�j�4������8;x���8)����Z�Y�]���A�Z��R��]FU����,�i`&@\~��!��:�ȼ�	vj��nr�s0���o(�y��Mr���GkZ�����7N��8�`x �x(6�9*G81��c��P[_����h�|:0�>'z�,A{��'���?��R�P]k�!+�+��NVFU�a<@d9g�D(�o�#�un�%��B0�n_���؉�ǚi��:�m k��w^�#$9`s"�:���lOP�����_.����r��Hp����+�m�zi�샏 ��/��1,�!��g�p�� �|%�3\�&����L��qׇ���N~4o#n���x�N`�I��U\�tv|��~vf�U��xA���k�'`ِ'��l�S��Z����;T֌L:����h�B�@$ؤ��o�.��0�@	�R3j��P�Od/�_�x}��I�I��}K��W�K��q~m" ��L�W�����;C	�2��ReIn�'Ė�g �5�V�kc��c��Xe�p��A�ښv�Uq�l����'������]��-�z�[��f����O2�[�4*��;��{��8�Q�o� �`����*<��H'�8�9O}��B��l�^T�,�Crް�u~Y����9���; �F���N'4Z���L��rS}m���R�=�]�)�V��ig�	ڎE�د$�鋡��{���@dJ:�֌�Ȼ�d����R�D�/!��~�&��JY�Ku��U��Py���#EJk�~���VQ�j+��@���1�:2�[޺7X�1�;]�56�=m}uZ�����n�Ii�'�7V, �k�y���~�8�遲C�f��w�1Aa���s�&�L�<���\1���	��<�������Y����xK�g�����c����}�Z;"މ�?{m�B�~��)z�>��0�C���2i�i�L�"��5S�_���a���i�Db�⮲˄��-�xiu�T`B#q�«=�#� �׫�(���tw&����l%o �C�Ri�0SG��b��v��Gis��@�g�Q�z��X<���
�	Q��%~�3xG��ϋ,���%����h�59���ņ�Y]�{N��[.d�Z�W�|����o���S|��.ƛ���4�m3�g�S�ԏ����{r`=�n�=+��"��O���.���}��\M���Z7I����7��.i�iO�Wp���2v�?j�5����`�ʱ��~_��$����BA�Q��,�V�{�Hƭ^j�~7o=��'>D�h�� �
4Hq��;�M�L��)��E�mE&��5�M�Zi�W8Բw�
�s#_+2��Q��a��}܋�[ѹ<�ͮ�\p3bk���)O$8b?��n&�sz��`|L؞vn�:8�5��C#��$�K'��&Ǧx̾��^�]U�=�e�i"�$���v�p&v��8��^�	��>U�����č#�W�	�vʺ�z�+���+�c�)�o�L
�;�`�����܈�,��j�߱�I��)V3/Zfw.z·@�q���M�mؓ+?��^#
�	z�.��vĖ�C����4 �R���nQf�s�@6������/�_����M�~<o��y�}�<�O��gV9�X$@�v$�AX�bp��	���'<g�=�����S�C�-k���n��tx��8m������^�.l�搣��}��m���}f`tT��П�y�3���u;my�O���2�x� $���XYٖ%3�|P��!�ln��}N��tj�<��������Wh�r�{3�ܮ��+�Z0���c��N1�y��%|�2�=-M�2�O��m�]S�g��T�>s�mu+�sOI�,F�m �Ʒy hL�?Xzz�p-1�[�!hA��Y��v�K^s����O��}
��d���B]����iŵNU�?�bw�NOZ��!���k�"�UA|��E���Y��%}�;��GZ���S'���:#�y7ϥ��?�p�6Q.`�{�!٤��}ih)��C=T]&�;���dYO�lևg�|�D�䃧��E�wx�嫔���fH���oNyd�(��}w��aPѿ���62��!�v��g�Y�p��ud��)&ښ6X�X���mLWA�yvx��]<Tݐ|Y1����z� 9���gl���/q�~Q����}�,��(��f2?�&�Ϻ;�w��~�����3@eS��p_[(Q�^8���DO�*�̀K
����2���7l���I�m]#0?��z`��A���*(��NS�U�
� G��3ví��Lq]�A���$k0��hCM�T\��^ �y���>�8�NP,�[g��~7��y��a�����Tb��N�t#�ƗOK�m�!�G�96L35�ze�6j��s���%��-x��BM����w�'���	�k��wq��(���=�.��[��s���ʝ����5�mB��A����&q� �ۅ��T�t��K5�w��H���%k�ȉ��n�h������` �Z��m�n�,z����fO�㹂'�ȕ��������Aə	j<ܽA"���x�#��w��e��O���_lD�|��x�c'O?FU�X�	���ȅ-��Mv��KM���S`������tZ��7-��ȉT�)����m��qB~,o0ᛔ�)zG�@��;^>�V�@��J�>�0�=�:Dg��@�m�_`U����f�>;8��rd����b�Y�L��{fN�ЩDoZ�
���7T2� ��'l��為
NFJ���]T�5V�{?տǇP�c�:o_��d��H7}߫]*�8.aO�P��kGV�df�b��gT�/�8Mc��g%M�&[�����)A���r���_L��1��)��
��0R<k�t�� PjB	.�݆�b�HW��aN8+� ��j K �u��3�4\O�`g����׵�q	A�u|gn-� ��Zǂ�J�t����#�.)�Ke!����%�Q���d�W�r��8����.���3�P��~_�^|���YV�ؼ�e��FzW��x� �vZ2�W(��ua�c���ЄFF ���ǵV�f���;d���ܞ�E�D�mO��0f��I! 󞾑��o���yZ��8���P�TgM�h�Op:3��6�s  �x�ҩ���3�*��"�7$r��k�����~�距R|@����=�fh����4�5s�m�+�Z�S��h�
@mxA��6d�/��ީ��IM �)nXB�F�����Mx�|]`"4��
0	{,�B�S%��F�K|q.#o��衳��<��^d�� �Q��B������-~@�r�+�Wn�m��6�c�6��l@<�l.���䝭^�󀑟�t������c��9���)� @�`��s�0�i���eޜ&썽�z����$�_B����^sv����	d,�x��V����p�=nq�~.&�gp1�+�p/�sic��pO�%��yM���8u���u0�I6f��p����B�{�����YIʐ�G.��!�o����`ZJMz�Jv��ÏøSP��G�g��?�s�;���S���>��^8~x��8��� +�����=��6v'����磖� �_��Y>��?��Z������Z�[�.�1ix�g�*"�zH����W7C�W��I�����@��Z�"<84�P��4��݈�E�2������A2{��^ԅ��װ�>�v�9+@Jw�*.��fl�[o�UT8�N��.�{��6(� 0�	d�Z�]�l'Ib ���i63�]���un���v� �"���n�h���xq��P�s��0��ztY��}&�S6ϯ��%�ل��H,"Ϛh@����[Izo�8�-�;�XJ�{c[P�[�<��=��i��n�Ω� ;�4���>!A	�;���%�B��{0��?�#L�6�t�o���5�=U5��q�����B� ir�n^5�b%�V�$����[ �!���#1m�$�����gX��s#�%��Xqb�e���A����_o�ג�N�U�-��n�k94�'O�T�s3T���XS���*|��Z���,/BY����=�[K4@���e�z���4�z�f7��%������!I�[�ٸP��7u��!�8B~k�Lz�􊶀m|�'�N��u�� g񠺠���F�,�{ۣj�M��O���k���b?��1��..+['0M�3�mo �ل����G(3z��w�U� ��l�ˀ/M�l-�)�iºֵ�ķ��.�i��f�������7b�RJ���N9���z@��4�˕y�n�|d�͘�WHߤc��G@��9���ς��y�\�9:8�u�f�#@BЌ�څ	=��Aԝ ��r�r�=�+q
�CN/�ʹǋ��c�o x�խ{mI��1D^��V6���w_Mi����0��Rڕ�Y��(��P��������V����T=����1Yn&R�X@-���%��Gf�Sq�" �J�"�I�+EmR�#6�|���� 
K	�J���)�H����F���˔4��n���i�xBD���8����ߣl��F3	����u3��`��q�f����٦4(y��?&ײ|zH�~iB��}���m%�[�u�@�LG	�=Γ�O�}o�7̝����kcb��Z"o���⢵<�MYz�|��쭔|�/ʨ�s�:<�-v�ÃQo���P�`0^�f���`�*B_I�=�',E�9�z<0��M�����~є��vʃ^�;]mQ%J���-׀8����0��◜`�R��g�����pTR7�!n��<z[��S;FJ3�kHL�$���7V0�P�ٴj�+
�K�F�厀_h?\E�+Vc;�	��OpE���9��ԣ�?	vG���`�)���X��:� ;�m��yؽ����8�]�K[���
�j<���ֶH���B1͵�/Qo�￢u|x^k�g
�k(<>��{����4�7���a�� � �K������` ��mm��e���5n4�(%\��ʡ!s��� ����3Y�N8��Zhs��F�I�ƻ탏L����u5���,{��9�!��M���w��#0��|8�\_�"a�H4./.f--V�\�,E�a*� ��wJD$k?��3��n��	�ϺS���	+�/��s�6�ǻ�Q� (p��O]�8��}8��Kh���*@����hΜ@\w��Ge�Nm����������^�h��J3�/����T3�Z���1����t~���#i'<�� ]�2^@�N�0aid�6��xO�#�����l�Q�Yl��dCS2<
r�9N�V~<��@��4�4
/�
n�P�D�dU-�8²��R���!�d�ջ�F(�zv��䌂1������plsJ��]&T���&��=��г(-��e8%כ��M��2�))���"R ��Ľs�\��jv�	�/�z�W�#����{|ʂ.��Ij�B#�h�ʲ��c�?��ݏ��I��_f��,~��� {fA1ֶ�k]{OqF�[�+�@�B���/7`l�k1<�ѓ�l�$7x6�2�FO��7�3�VZFx�����K}���?�69U��'vx$v�y?w�9��5��_�Xݽ�]N�����ĸ�(�������~\ �i�|%ĸ���m�S�A$�����ń{lsY��{R���K��{)a@�t�9���%rk���,�g�au|)F��'�x�nr�|�g%�����vEl���~��(=�
w�s�)#��|�	�������?8� �q�š���,�L{z�}��K�z����w��˺�|8�_��s� 4>����L���[��Hu��n�x��w�N�K�F���G�fj�\�2fzU�f/wo��K����G�&U^��f���F�FWS��G����\%�wWv��O�g�O��,e��3����u�Q�>�y��u��Q���J�����l�Y'�6.�VQ iS�;���`LZ��Jm�EZ�>�BM�����V��UO��ۣ̐Lξʦ�/d�I����-ԃ���|BT,��;RU��X�N���[���˲J0_\���m�-[v.���R���Jf�����fi�	 q�*��<�C�����Fn�O�B����Dy�Ûog�M�"�B�:���D�B��o���>CN	"�{Z9cC��<}w<����M�����Y�̓Y�l*3�8��ޫ�J���Q�Df�1�e{��_ޟ�����۹�u]������u�B��,I�;�����F�=[,{d2t�-S5-1������+@����(9��!Jk��V	�K���{yh:��&�����1aZd��/C˦~T��sv7�M#�au�^��2kr�Ej9�'�G>���*S�-*�_�"�+�*񐳷���w��A��|<��b� �պ�y����~��r���؏��웅��Kr��r�}I���ȇx�����ś�j�wh��k,J���(�����|`�P���}\�R�m������^���s\����( 9X����@�m�}��y���n�\J���z����K��n�9��Y�FV��@JnP�=X9�Eʐ9b��v�5���`6iYϏi�R�^��**�ܟ2L�a���7Y[� J��kρ�a:!��2���Y����<�~�{p�0;�9��h�
�%܄>d�>AӋ��ɯԑ�jD2�q�7Z��ݟ��>Xe����[#�Y7�?z�y�]*	�Q�
L��xGP�͈�I�-wX���a�ʱ�	��Nc�yjl��F��U>��=�:��B����
gN@z��K��
s��X�VH(��],���:%=#L�VW�:7���dߞ�Q�?�F>D�	�~\����^<I�-��n�Q����6O��;9|��"��%�}J��=�:������	���d�Y�9�f�#�9�"� �6-, �bp��7�c¸��~D�򼷌�U�?��KC��c4����S���?�8="�g�	����'W��r��1��@��^�g��S�����v�-���o�/왮I�lؚm�G.���[���C�̷�v2,Lo�|�o�3����g�V?�^_��b���zX#��t����xK��aMy�����cN�W�K!ϙ͌�`l貘N��TM�r�f��\*��4��."ԥt����j��`�&�i��Iw�����ۻ�?�ȌR�Ro������mǅz��]�s�:=O�9�x�LVn�C����E�Н*:�F�#\;�2���u��;�Za^��yr�Cv$�֣܆S7E�]�ݲ�6��0��|�@�T1��F-Y�;��bb�u�-&�<����\Zj/�� �٠�D�M��~F1�� �����N�-��ۨo����ͮ����0B��{:
Gs��f��E���v���a��i���&�zg�
7��D#��%��)٭ȍ`01m�7_ş��r@��pr{?�_l�U#S{�� ��2�Q���S�h��_&��#Ӏ ��zc?� 8W�E���
C���2��8홲����2O��qyn"��=�.Uйg�.�sp �Q��D�f1n�MR�x�[�oZ��n������r
#����N+�k�H	晡���ʱ�U�I����8�2ۑ�7B~�~TڞFZ�b����EF���f�@��+��h�-�f���_�ؿ�O9�[��i�oJ`O�B��,5����76c�V�o�޸����Ai4iP���  �x���S��a��HG�6(9�Ӈп0��*P�a����]��r���wJ�_.�؃f�$��Um�Ko�,�b���X�9Q�|���tnC��v��OL���j��3*��
�gŕ-�SSYE-5�'B��Z��K��0� �é��r�]��O$�������3ůTc
�nӰ�����}C�	�{)B^�:��c����C^8�撆����΄�pc��ra�+0��Ϋ�&��c�sPhac�=gK|�d�N�9�4�̡�Ղ�~�Ey�M����&������W��1�|���KAJ����p��z/~}�����'v�i�қn%/��a��q{v�7%��a���}� �x+iu��Jw��/�쇞���E"��쵫��8��M��MF�YF�M�=��z���l?x�k���Ԙa��M�^T���@	�r�=]�a[l3�3��i��e�vp���A���m�x�г�C镧���J9D.�Y��9�=�����6�d�6��(�Ѝ��3Y�e��@�G%W�f�/�[�HYЇ"\��5��>5��*�Q�9$�(��S?���A�S�mqkڞ���U��_h��m��U#<���^��d�����@���pz3	n�Й��.}n��F��|�W�Z�s�j/����� 0ջ?��U�K�&��W4��qr�K��=�M1Խ�D_ZM����m��O->�����{�~VG�o.@���Y�z�ˠ;,��u`�S�WI��㨮�7��@�8鋡��B�� �٨�ڒZJ7w��/Ԓ&��x�Y�u �Raa���i9}Q��	3�?�B+��R?5=�=:\B����uҜ�_�wu*�����;��Q�N͔���(�P���ٸ��P8�k$���䰹�G j�Z�;)# T�y�[?�n1�ĭ�MbV���cD0��|�6g��P
d9s/֖��=Q����G�S�!��S��ײܛ`��H7/���n����~TaQ��P��6����1�?���7Y=��1N�S��Lob)Z�M6vv��4��Q�Z޼V-�0	&5�#�v��Z��,�Onn��i����e%��2�΢�r�'57aϠ}�Y.�{�^/��y�ׯ�D�u��|LJ���9�T���ڢ{���'8���y�-��^�,�	t�J�f��ۘ6W ��^.��}(��t=0�8"Oo�Ŭπ+�3=w#g�g�ޭ�B�}�������-J~�3dgl�R���щ�'�w�(Ãgq��:���0)��M����_iA�܉���|Q�P��p��hh��r<@��UN�H���&���q^���\�'�te��韱�Aī�9�����&�^Ka;Mdr�}���Z�R��q�z��w�Ȃ|1�!� ��'܀%ƴ�π3��b;��*��|����e��SzX;�i�rf�0�&�ɚ�E͍��]4�$�����.�C������3�T�D��~~�T&�%as7A�~W���κI��w:�^�����e�$z�2�y�J��ZW>Kj��<Q�;9�̿C�[�_P璍$�y� t��=?U�A���@.�0C�������m�5k=��:�G�!C�M�!��9Ps�R����_wZ����ǃ�`�.Q��)F�Ι�¶j #J��DAG��7��=�Q#Y�ѹ���2
\����H+�-슥HK��S�c0?S�K2��F(�S�N�{5�D�N^]�F��4��6^u��zߩYo�U,X��n��s�O��!xN���`�V��}�	���'.t�l� ��;�=��$�%q�870 ���E�a:�fP���fƀ�KԌ�lC2}���-�s)�/"�f�l�O�@�m��\F;]Z�m1�;ɐI�c���x����v�UR���x��Y��j���62ŭ==��� �����9��1~��^C��7%���˘ռ�]6�����/W��ʄ�u|x�$ҫ�݌_����P%�x�o}��h�%��Jٺe���}�.=@B?X݆-��7�O=!g+���)�<3x��%�Q��{��ҁ�#}j�H�K�uu
G*��(�����$[�Q��/��7\�W�1Y4��#��#���^R;^��o-U<1%!��"�F�x��M46�3�с�΋��N�!�n��Q�U;
��ވ��Ҵ{as�ڪ����ڳ�AH5�M�;��:�	��^���Zmg�.hCG�h�!�GS���4Q��*�ڿ/q�t�<�A��3��#;�������-�@=xw�LK+j��!�)�N�R�_k��oy_+��`.f�w@^{ω��h�R�
e "�?��UId3�e�n�P��Go4|4x&�{���T�^k�}������56Ĉ�����D��jy;�:wO��>�&�ġ���"�Sp&s��B�q�CS�s<�s2��*Q���j(��h��G̣؟i�Q��;��{o�Q7��r)�?��j�Y"��~����2���"񲤋�b��3����y �i�Β��A��2b���/�;,��m����-5�ߥ3m��H~ŝ��|+�J�AfP^�g�is�~&��9=XO2��$���vʡ7U�<O��� ߟ�.�H���9�� #;*I�W=�����W���2��o@_Ӌ���S,3]T���L��*@5���2m���b8paCq�{���i�i�����srȒ�|�.�[n?R���o����b)=�܁�"�%m� +B5�Đ�O����&�:�_���F޼���x����^�vw\��ҏv4�<�ų��6H���r���	��>i�4o��Oe����%~��F>�MZoDg`bI��e)Y��kl� ��@�s��^/���҆p�0@�Ac�E,�X	��FiZ� ��s@�[���!�Z}�sT���?uGZx@�פ��)_�?|`��G�s���:p�9�6�����S��{�@$U'{�,�1�����l-�z��xl&3~��������/_E"�9Hu���W�]�BZv� =#����t�掦Cıϗ�T
k&bt�@��ӭ��y������4y���lG������r�,$Y���lٛhBˌ>*�GK�����.�#�[�&tx5��V�4�ٺ�鏬���`f�a��48�'�v��۫�׾�2{I��Jt$����Ķ�k��(���_&���	O&>"�#[{�%D�J�)]c�n���&�N�j:����	U��|N��W���K��f6���K�)0%���
=��:K[B�W��Sh���f�}R�ʌنsk٤�ғ�W�G���M[憸O�Þ�{��nu߹'��Z%Di�1��cⲟ��|�V�~	���B���/�6�j&i�W��ȣZS㙿8��؛n�K��J7�otCF�{Gx78 
��냑�_��⽁��+�K:�[D{96���B�uZ�߆�NCי���r�q��i
)�B7��KRy_K��v���k�0H������j�\2���4�0�iW��`�Nm����
���%��j�(�KT?+`$"l�!1��	�,hB���w��p-c�h{����[��ju�8�'������f�0��������Gj��?����eb��!�%��#y�sb�&M�X��y �{��
4�p��G@OC�I#�8</����t���Q}��(�aex3s�¼�̵���P3�fA��G���bݻ»g��}yyH���/�h�M���[]�+�]�X�k������v��K/!A�*�8�!V)��l��F��)���Y劶,LZ�0t��y��y}��l�����@�>�M��� �c�hE��c�����J>+t��x��/;J�ZK~�!�xaV�Nj���{юXɚl�A�~������G*c�Qo���( �C�`�qq^'V�z w0f��X�T��e�H&��-u�'d��r���ܵ�I��	�ݼ�}=����J��D�1t=)1�D).�1�Et�*]X�7�/ԥM.�4��IS�K� �{IԤB~�Oĸ<��k��* �醛�xL����!4�qR��=��\tO��`���GQ�� z������Ҁ1x�X�j\��j�?t)��N�J)W�eCɓ�8N3��l��r��u2���uy���Ⴧyz�+�5"l�f�"�/�~>���;�jZt�^����,�Bu�A{(��- �_��7_ķ?V�g�T�?�p�C�6`qs��V5b�i�(ؖ�	�V�AK��OUu�_��o����Y}	O�)�C�;����>�ދ>-Ln�9g[�A�=����P�g�����H�g,�z`}���5?: �gU�	*n�g���4�ź���������@(/QRם��k�#;-��^��o;�4�mvC8k�ø��x���h2'��hp�G�ui� ��8S97�-�����=�d��2'�?a�:�h��cX�lT_�n��o_�P���Z~��Ѫ�*��yX0�Ɉ�|��������xQl����-fx
?(�\� ӴG��0}�����M��b�T%�+9RhΆH`��ߟdb�&z�<\�jVN]VÒ��J���W	�dq0?i�u�r�a�/;a�,�$�~��A��P��@�N��F�O?��j�����a��e��J�������I�33�<�*$�ή\�����7��p��T� �[�D�/_�
Gג�-�ɀ~�����z�+�Ѐ%��Xek��������y��5���G�)��;��4g/��zF�F'���%��L�/�h���<Z���'(}�mh�e�,ld�]5�F��-����u�Z���t�~K/�i�_��繹ͬN�����0�]�_��:���X���>t��?"��8o�~�Ys�䳫�Γ�Z�q�z�2�T�1xXA� ���(3�.בe�b��My�<����u�*��Z�Nk��9�vۅtl���af�����������bC/�̀$�R���)�m��llCs�����'������	��ȶR��{��[�*��P/��Á����E����ewP	���n����w��<�B~��@DL�J�`h�!���XP��e�Tȿ��rQe�s��^�19�����1���������=j�cC�u�닼d���b��YZ��t]�o�Z��^bY#*�W�-f|]U>���]���^>�֥9��Ѐ�wh����E�͒,����d!���qexSR��v�;$R�l��������*���4��v�/O���3�V2�#r�>X�D�#@Lu�T��4G9�,�����4`� eP]Gjn�o@�\1s�>��3̇X��9�#���`̓��X�`��ћv�?|����_����	vC��~Y	��#�.��ri�C�
�.%����>�%�`���_&�|�|榀����|��ptʕ���Ȫ-�˙��V�2��:r�^�xt��b!�7=���0v�2��P�F�(�3I�<,r���g�o��o0q����1����v�q��r�E>�C'=����4G�f�����&���7��M?'`JPRɖ;c�!�_X��T7���wO��WD��Lh�w)�oC1��m�������6��@s"�IM����}���Fq�O�n��O�k}Qx�V%���B8M�d���2~D���2�2W����>7�叒Z� �&���V5�N?R6	<�F��Ke�e��6%J�&oX{�������?���8*���l��l 1d���y!����!-�)�s~�8���G��'[���S��'��G�^���S
�����4�r"	�^���<�q�*�0�v��8���T�
�k���(�>ot�+^�ry�h�ٜ6��q�m��t33D:)�1I�����)�����ܑ<��Nw:�x��k���Iʺ���)5�>q驈v�����p�g��r�R �A��O*5m�Y���V�B��D��D���M��G������b��������D�����)�R$�:�E���j��@��2�D�l�ATl��@ ����M'S�,��JUj��բA��;�p�HZ�۔�X���ڷ܎�>gA� �I>�תnH2��0�!he�����<:�ʥjW������so��~��%�A�ݎ����D]3�H�6S�荗k�gV���Ȃ)�{�0���l��sv;3R�k�D%+�.�E����I�ŻILNK���%X���{�T���̠V��J�9(� ���;	�����F��-T���cL�����N#�1xs4��>6�-����}�PU ~�T�	����
~�TZx@y� i�勧t�黎��?�F���޼m�����4��L�7�)i|���ޟ���9�q��cC��q�|���w[lR;C��7Q��E;\�]���R��|����\���E�P!����T��?܅�Mw��;G�D	��^���`�Xj&F<0hb�Dy^�@�p�B�����^��Y�vD+r�Nx�t̠S�r���A�����愎WW��>K�pIX16o<ͨ��MC�V ��,�� Խ ���jv34�d��)`�r���oz�����^�gf����W�dn]rf�_g�J�?�1��Pj`JAwE�A8��Z��\d���Q��7�L ��F�Y�&|��V��-%S4>�ZJ�h��c�ݨ�VY(м}Zt���J%Q�������-���P�Ə���<հ��ws�D���>�~W��GQȞ�\՚���?@������)��� �abdy��m2;�1 �t�oM/�AԈ^�;G�.�����H�J�e+ɔN��y?G���>�+�;�]�j��|Ql�>�����dg:~�(`+ M�����<�Wlb�.���c�>}R湾�6�B�vw����q����e�����j��pk(*E`��曣3+��tI��9A5��R��J�*"�����;2sZ�a]��/�}�sfR�z4�'��?���/�o�I�/����X�"���Õ�ڴ�|gL�Z7�o��?�a�w�9�C̞���~�I����M�$�����t̉��Ǯ?�d�ٛᣛ�*�Y�e�QB��2*�5��ח6O���.�}|����įq�G������!��O�6ة���i��d�� b%R�=�J:��4�!��E��\*�R�C��cd:���<���O��1�����!bz዗�j����]i�ii\�&��vv�r<v�#n��ӏ��i�l:Տ6�+�>&4Y�i��6�^���ۛ��
�"ݯ�]�Z/������J�/����G8�z����q��/�\e5�.�&���b-��l/�l0�8)q9�	ṒH�K�w�̤[��_�	��9�Aʚ��8�� �U��4Y����u}�S��3�������+5�yf^,$�����bކ��Y�+���ۚ�y��f�gI�'�ӧ)�M%�6M�.-�ҕ2����{Dac�<�;�HUM�W}�v�����|Qt����ǿ���$��l�f��}#�'c�X��OX����L�ѪU��<��f�$S�h^z�L�B�W���#9�6tnӵ�4�"�砃G�'VW��O���`}�<n�p3X	M�J��>�뜃��~�_����gX�8���QV�Cc'�=�?��
6v�J�5,�d�>n�
�UBJ�riMw�����W7��;��� �\щN]bљ�{*��A������hZ0~��&%�o����r6�����'ס" �w�g���0�s�ׁ��˟� �q�jz%Ȉ)�w���/�*�#H�yϣ���~k�3i�SlE�
)���'�xO6���.'t^$�*�x������`�Z�2�)�L�!�7�7�<H�Ø(�2�Qn��,�'�����6M�kɢb�VX[t}$&��E�̫�EB���d�{(Mk�D{�Щk8%[r�.voe5��t�R꿨�?�K�o���~�����V�j��6R����zT�h˶26��ל��8�c덈xDV�],y:ق`��9��{#���tV�T畝�_VE@3�{�ב5{�r'�X����=�"�N�;���N��@��<g��;0���J2��-��fC��D����ms�|7�;-��6,����>�Ǣ�C��uW47���5R�����:}��il��y*X]��m�F����~&����7Ȗq�f��I�?'W;�v��FHN�_#w�r�S�����"
�-'��yy������ ��Oi-�vG��}�J:�&C��#|/��_-�U��z���O�z~H�7�9y�B�L��������%Q�X^~�cy�\۞�|Q�����bP�5�.�#�=j�^}�*��vhD�Ə��eo./�[^|��Å��99�_�[��C+�����>�H��I����r(;$�w,/�6������Z���6��;���$;;?a��T#��fԇe��_�p��@p��eNK���o므�f�dd��;��ڂ�ֆ58Y����Ϩ����VE��:�!��_D�"�8]��x�a��+�C�<V��?��J��$���ze"��3����^�f�0���~G\"f	�,�%v�y���>���͙�t��+s!�Ƥ��osA�������a4�f%��rl���lۿ%\��(Y�=��[w_٢j~[|�}Y��[�5L�r�BhA���"��]b��C�/u�9a��$պ�z 
jy���ϡS3)��
�:��j�8�b�9��S�[�)��J����Oˋ���w}?�ހ���N qہ�ݧ�%�S���v�L?������`H`��g��4�C�ץ��N�d�Y62����N��Ԑ�3t��P�K8���t-�ic��&�t�)*��Z3ٗ@C�=��5����}��ӗD���.�
��'��Jտ�=b��|Ԃ��� 6 ʣ��\Gŷ�j)y	IϞ�%�
���yQ?�cv�����̵cA�@�?,����`|�M�8���d4���i������\�ڵ����H����j"\�Rl��^C%b\�ea��������$LQ�KֱS:Q��Y+�o�Nf�0��R@/����;��V����|��|VJ $��1{�3%�6�7�BO���-�Y��U3�FM8<	#���P��NA�=�1�<��V�*b1Z2���_ŝ_��1�Y݆�|HK��NJ�'M��s�fo��tn9�Q���c��3ÕP���_!Kjn�fw��vz7�j���١�\u�H]:��_��?hy)�=E���>cP��6�� �:��eM8^D6�y��?��+�vo�GwÛ H���G]��L1�R1*9��q;K&̕��p�v��ֆ呉�����;f���c��a�[�Ė	[�`4G~Ɋb.�Q�d(�N��L��#`u;p�l���HWR\�b7�̬�L(j)C�ɬ����P᫪08J y;�(a0���׹iz�(��%R/bP���S6�B�� �[�~f���n@7���3����Aɟo����<&6�}��������B�t&���h/x��Qq�&,�C�v��;m�s���I_��=`֎f�<���d���sc�q�VH�w�}Y}�/:2r�׬*���y{4�!n�G�{�����4ۤ©s�hG`�����\S���E�cYKk�hθ�i�_�	!�a^.x��v�EF��2Rw��~�'�������D�CL<#�FqD.=8��|�v��}X̅t��11S���J�fk5>����Y_M1$�'I�s�;f���w�;��❯=~��A�1ߓ� nF�y�ۚPfamM���!z5.��p�7c�5C%���4��z�h�M*C��0oOK���Ǡ�+~��&��˫*��nk��٭)�Ei; ��P]����z�B�R<���I0�٣�����K�Ǩ��\�CN�>ۿ���/�2���=n'�^)qym�ក�S�����'J��-5��w�F���{8;�.�l���ʑ#�#�1O��]�z�j)�8�5���%4&��ݐͯ���ܗ�7��k���p|�G��q�]]��q�+v���gV�i �/��+��R�HUg�p�e�Ҽ��ο��J������R�Nٔ7���BG]����z��� E��p9ٳ;K�<�ݼ 92r�}�Ϯj�&�!�U
N��y�L|/�L�s0)�Jx�ͯD0�,�V�����
���P�ɗ�B���̄J�O�G��G̛n��Ij��R�l!��]O�R$�\uëJ���Y�uO���j�bN~, tX���H���/��ĩM�?7��q�,e6��l�R9�e~��
ɑ��]k䚴� U����_��,���77�Bx�ڄ�w��q�� M������.�!/"��b�)$�/��«�����^
��:㌝K���g��M���e��?Gީ�J*��vJᝄ�٠3J�t���Sǚ�3����̽�&CbKLO����jŅy�|ؐ�Z!��0$m2�^7�a̽�8I���5�b��N�Y���TJ�FL{���a�dR�#ۋ�9R��Au�������,��	��WL�b�:3<�����'}o���b�Н�~���c�L�q��
���a=���M���9-����H�Lyw���;I���\kvD�Bz�Pw��><�\��`�Vg��}��w���Y� ����^�ݚ�f�j��(����gC�^���L��EgЇ��9B���ܓV\c�F#�4�����	��z!�f;Ԓ��>+{���Ӽ��,9��y�f\��[�,��)�P�	�V�9L2��G�>n^z3������iV�8�l�Q�NZ������I]usώe��\i����w���	�b��/V�v�tY_iB�����,��{�z�8�Q��۔�ɏ�1�g�
8m��8�2{M���*^���2:EC
0��NG�H�'Gï�sE�Tf�f���l��;:���t����w�pH%�1N|�җ�=S����&1�@�����9E����-���7���!�][�����q�dKL�^'����Zzjo�|�7D��!r��yU����9�ӊ>���WT"h���f���!x�C��$�Cٳ�e��g�7���	ϝ������O#]}B:w(����Bi���V	����W�j`
��l�ī����A�ES�ē�FN���{�zX;y/&��dpJ�����Nj���n��Q��ߧ����@�Ik�a��>�Wei������h��U?C��5+���ƻyP��8z��F~��k�v����#��׶�6���Y&dz�{�7�ǵ�ԭ_���y�{ډ�6�]x%AÎ��d�wO��to2.�(/��q;�[d@�i�nةʜ����m�I�P�Mi�T$a��m�)�E���7q��c����KrO��=�+*StPr�{zȉ��<�=��t;9r��\���CìY����tO��S~�^�_5�c@�$ua�oh�����7!��6n �fG��ﲊ��3LGn������F>������R[U������U	_���@:�\V����n	��=k�&*kGF$�~S��|��q���GR�)�2����i�:��t�&��d�JOTVo��֞�������Q���'���Ƃ����2/���� ��+>�v2�K� W�X�fײ�9{�52����R}��}U5o������*4v�F��\�wl���]���\���t\,E�+�ݡ�D�K��z��&��^�s�E[���X��jZ�ѷKݠ[�_T�8�_�$�4��yL����B�W�h���W�Ks�m�ַ\��8�A�ǀ�t����iݲ��slV�z�k�`Џ��b~,cV�$�珖���or�/*���Xi�r�}���W-%��˿?�/C�G�e�A������(Y�2�m �k����<��'���~!�O�@�8����W
�z0}�����\�/�ۓ���+?�g�3�X��/3��y�:C����[�>>R���uc�>;�h&O�_�	,���]�o��c��Ʊ���	�Wo '��-��*�^x�9�f��Ǆ��v��z�R|I^-Y�C��U��ɣ�z]�M�cP���kKʡ�G�C��3s:T�f<�w���m�dS6ec���ԓ�I��������w�7�>'C�������Z6�E���ݢ�ĕ҇� ��*<S�!�����������.��ǐ�]77\��o&1�Y��zOI�0�{2"��gY�Ƴ.��it��ǐ=����6��3�l��Ǘ-	4` 61�A�H!=*��I�g�X��P�Ѣ:���|(��уj%�����T�OT�A:`�W�+7����7�H�iR�<��]�:�.�Z��ؓ�^p���,����$X�p�jᡌ���M�u���noH�UM�B�H���>��6��YI����[zy���igy�Ŏ#��8i����"P���ŗ�{J�����	X1D���xM��
��L�����iUw��8C:P�z���R�^�h�gh[.��$��0W�F��|ȗ�������NrEE�K}R�'�V��
��o6c=���Bt�C�L�8�c����8�,\�E�ms����|��f�v�V ������w1�6s����0���ԃ3muR��]"��	���x�/�9��X�]�"#���P c%>Pϧ�"(uUQ���K-f�����9��y�SBsaF�a]bN}6d0Z�$	��(�X��n�gn.�R��-�ň�{��a��,b�6�q+C����F�.(x�|������hޫ�{�ǆO�}��`�(oIn��,ύ���(�fւ���,�ۂ��(�>�9�����1�a�U^��W�1��<{�x�ttYQ��V��S_�K����Ճ�IJo5R�m�𿊻$�
��o��ҠI�����D�@u�2$'�W>:� ��"���<�02��Ne�Ɣ��dǱR�:hB�Ʉg��g�5���1ֺ�i`�����M��S���"�ܫ��,2v)Hܪ���~'�>\=CM��s{G3︌��=�2�b�a�̙�nŭNx��*~��Ϣ�撪���	��v��w/U�ţ,RNT�chI�+8���m>�]��@��v��EE 9ʰ����L��ha��Q�8�E����i�݅�Z����Z�jE-��j��J YU�YT�f<9���۾K&5�ýU5����l(��#I��ɿ�x(�=pl����2m��F!��'������f���������DA$�=�1��Cɮ���J���z�����O�W^s�Ո;�R��P�����l�襟m;ʝ+��\��dr�&la7+���R��Wv��^�5Tv��5Ѵb��'_���ܕ`<�0Y��H|����«�f��	�W	�oJ�<�|��j��x�';��Ɍ3��&T�<W�u�)��� E��owP�y%@Lj) *��M��$�k�/e������U��Q'{]f|#Y��z噺��<�o�C���2���@��9%����ަ����\�Ί%�p�K�S&}�5I�19O�rfd�lrp�7$�PR�#��:XN�S��ss�*gk�ȥB�W�e�ڱ�}�4o|aq/�� ����-X#��g��փ$Ǹ�YV�H{	ɟ�d�> ��ǎ��1�b��`���������c�r����E)"I��C�����6�_���l�Mr
�P���`��ξ��ǿg��Q��>��ʢ����Q�?�`RoA/�/
C
&���_q+n�/���~�U���İu�R�Ɓfn���,5��h�y�R_n5�ڳ�`g�vm�|]�U8��8�9/�9��|�>�	&�t��� ���f6�����>�{]P�z�h��x�{dA|p����=�%By�&`��2��(�ab	���3Za#RGeW�D�x�ـ��Z�j�{s%�~.�W��~^�b¤�G����#!��O�ZI]x#�k����j���rP6�T�:������{�BMR���ƛ�l����k��J L���
�_�����vxQ�~0�ݻ�y��/"<N�ۧ!J�d0U��ךy�+�&��r��o��@o|�Xl}��$8?��j9�s���O����)՟�@?7j��!�Nqf5��[��h�j@b���Bc�K�NGa��H/��G�h�P�t�:�7E��K�V:�y���_*�c2�1��Ll\�ۨ ������4�IQ���dϮV���v��)����g߀0�1�ވ�r�t�ฑk/��M���o�ұ�c5Mg�վC����= ��Q��)���{��\)�k'����`��]XP��ի�i��3�V�-Ѹ�;0lm)��*�H�b��K!`]@���)Y����z�����c��Hz��={�7�*���/o�z��ȝX1���B�,Th,.)�)z�١Ѓ����~�|�l�JR`tQ M?��L�dgǮ�`�Ȣ&P�H�}wC.ab������{�|�&T�:���N��a�#c�i�^Y�J����{�U{���U�Ʉk�d_,#��ۼ���˩51들��]����Ң����W�������+�!�qk�S@��w�2�J�!���;P$.Q�idI,�][���ah|�7sNol<ď�}��B|����̎�Nu���kZ���읜�﷢�A�:�tYb[b�8�7UH�_�����;�`kd�X`\�<�`C^?�;Z�A���}��=��BDyQy��sGc?�b�l4�p��Z�z��k�EAV��6���:w��[�o�;릧Yt��Mm��w�v�߄t�����������JU�O����0�PA,y#1�?����7�E\�,�$�\#���nN:/�y���,�g�z��m���̍�l'���+�,�f��������� L$�$�6۟!)�����pm6{��������S'�����jjSK����WWd'�=A�_�f�3���2ԝB�ۖ��a�W�k�Ò�C)�b_&:'�0&jF�m�es�B��SK�����k��ƟFk��r���|�C��R�A~�]F�f�=Ce�7>��1%�e��%3�!ͯ��۸������Xw���A�K���@���$�k v=P������a�@���젬�:�Ȥ��z^��'�����H�	��޽�^�K
d�1"�Vy�k;�G�d����l�B0����8��4D)�`��ɟݫV��|��}]%Gy�̇9h�e����OM�;��wnA7E$S�A�P�W3��t���I��v�z�����f����̢�:k��	<�wK�H��Ԥ������)��Izf^�S]s#FPޤ�T{��ͣ&���t����akg!r~�q���ۍ��G�&���1��Q�Sf��d���`Y�IeշKG|4�5���@O(�(�GI,�h��f�!5�i7����T3����HA����!�i�ϯ�v�56I�Q4���KP�m��or�Ъ�ұ�ď�y_mw�^�6�
k��	�D���&�ҭxb��)�3'o�������5���PK�ho�ipC���羄U�:=B{�L$����ɭ8���c3v�7��q�r�s���c���c=�����--����0w��x4_^��|�BB�Tq�ޙ61��{.(5���Z^C#dqw�ܑ X;�F�&��.OXC=+Z�qj�"MZ#7h��&i�w<0c���cB���q77��Ύ�(����4�~�^F
�t��\g4�`Q�2���v/N#L�7�}��\�G��Fx����;�+�T)ʙ==�?r��_X����`���k�%>�,��|�2{R����iQ������M�]�y��z��D��vvef���榒7V߄�=���\��`?Sb���#/oN���ȂY��;GE7�Wi,IW#��MwO�a��b���ޚ��|�םx;~�	p������������=_��H��L}V�o|�q�e����ŵ)X)�k/V��<���#�/�s0�Jd���S�~�,�*,�V�x/�c4��O)@K�Qx�ry&P��E|��Oo_:�)�����2,�.jF�;�ARBi�n�E�����pD�J�DA:$Dr �.����w_x?���y�~�7��ڱ�:�y����C�qY��<��Ji�(4����g���?o�ѧ�sZ�G���j�P���{бz�q�����
�_A�p��\e�N�~�J��t�AC�I7�sZ��:�3�"$�oD8�^[V����~0h\,�,������2VgV>a���p���ŏq��>/[s�4��aW�M]��Ǐ��!Wg ��䜴�##9Pѭ8"&ذ#�T�c^���\�v��]����#Z7U����^�>�C=��¸��T"r��q�օ���3B$�����E~���+�>����iU�
�ʑ��|A˪�	�׳T_���m�Y���91�����a��]3�R}�)�U�(��/���ױb{Z�����uJ
��k��CZ���/َ[ Py�\�~Ԛ��|�n%M⩕BeDZ�c�Y<��7�e��R�&z��|�p:U�Y�� '���x�/�Ԕ�f5O�-ef�~sƈ�s�X
���Y���U0���/�{E��32ů�]���4��e�I_�%�X��Lf�iXy���1�i����}<f3�|j���I���ʫbR��������%�_��V0�|j _I�r���nd������^i�ZM�>܆q/�,��]\Li�'��!༵��Ǐ+&[�cʛ�l>'.�Ӯ�W�Qvs�6�.wTF4�(�~�<r݊�g-11H�Ͼ������sPy N,�����/�
Z��\ӽ��n7�q���Vڙ��kY|�?�-��1��x����T(	Ж,Ws�Q�Q�*��9A��P��;�b��[6'&�������Ql�r��;���:��ǿय़�P�2��A]���'g��G�7?���
�~}�g�aʏ��L�q����g#f�������(\�'t}a���.����$����Y�×��Pd?%Ge�$l�E�G�h�Bި�X��@u�r#��2\�y���T�|i�!�K�sN��YU�1k;�uTa�Hn�#�]��N�~1q�I��m��_/.�>��,e+q�"f��9�ϸ7�CF���*�2G=���������'v$WoD�v��}�I�y�Q��� +�4g`E�����X���ǣ����"��U�z#".NB��湏7���T��no=(,�\�J���dW[���WTQ�b��X���٣�����W�,S���������D�l
��������$P ��=?~�.���u�R�l�Q�3��&�T���T	/�`�b��/��������·E�׫a38��j^&��Ud/��u���&�ڊ�b�͜��y�1�頪�����	��ɕs��v8������'hs�7���Z�:V�����o�� se�`|�6H��C;�v�h:sv{�	��\b~�iҪ0��L&2�_��X�*�7�?�ַۨ��#�<�1i�q		���k龬UM(�槑㯿$�'m%�H��h�"p<s`Q�lQ_݀ZkZ�ft����H�&uH��9^�H��^+���>���u��_��P�ݎA'��᳭�5�/��k"���b
{Ե}_~!����`FS!��\b�g�AMg�i���R^Wù#��I�U{Ԧ;l��-��a�^�`��3b�R��\Yv�jL��N�u5S�DB���.M�|���&�\��[��5�v�-�G���Y� �%�&��0%�F1���-]��V�?"���S_��lr_dڗ�.qtAz�)0�co�Yڶ΋��m�	rS*[�й�yV`:��0ުd\ �@O��|��$>�7�Y�؆�lL$\,0�r�z�{V����e8d5v0���.�&M�����m->ַ��Mn�{`���)F0:|��T^.��m.����Ɨ�kڏ:6�f?W �E��hM��sK�*C�����G{+�g�$�I�Q�$�ɵ-XΈ�H��r.�繆����P�""/=��C�����#��;{�+R��^��U��mv���f����g{���� u5��<��Ą� ��h%��� b��=�Qy�D'�o�<k��W�-&�z�	ɏ��ր��`v�p$�$�k:�"�U�: )��I&M�m	's̖dRy��2�sf��o׿���P9oW���P��yU�}|_hR�\����JAh��Lx��b5$�WNm��|������Z����������o�W1�:�~q�r@�3-�L|/x�D;�Œ�����y�����*{�v�{/�%_e��G`g�����Mwj�ۏ��L\��*A�{N䕞���'�����7�K��]�@·�K�nނ�1x��'Šk��_���[s)c�ڍ���{,7v���8����)�9��`C�&u/x�����ވ�n�<��)HIP�*��cZj'1�Ռ��C�q!����8!�|��Q  ?�z�ޚJ�ԋ6���M
��H�8ѯ��&-g�C�>���p�?�
ǣ��5�:��)�1��GEQga��H"�ą��
>�XE���!�f5/���N>|�	��Ԋ�/��M���	T�����E��H�5J�J\�U�����_�ܚ#��;\�T���M"
M�.��B8���o�3���=�FYͯ_���,�4m�^c�!˶��F��qB�-�uS����b��������ҍgm��Jc����Dq.��.K3��hմ��퇅Oy̓Y�h��(��Z)���1�+��Hez�ě`��*��#���E�x�t��*t$�������-�/�iՄ�;wo�_��
PrkY?~Q�i�_#�lhG��!@��� ��-�&!e��n}4��$8	A��i�B���dp��wWSx�#��nt��ֵ�o�cp.�/�ȓ[��M�MhO��;˭ ��U� p8���S�~ͫ�G�����A��/�Zwb�jg���G%�Ŀq���J`h�sA)��Y�\�����%N��1��n�.6&���=Q��m]���������(����Ш0�Fv�~��jj�X cy��ҵ���Hs�U��m�8�YY�މY����1�J�
��"�gd`rʟ���Մ<�Aoj�o�4������~͇�b���T���N�9dZ�����-S�<�5�AX�|f<���a�������~�Lb]C/�j�����f"� x��{������4	u����_�0�͕2� ��\�m�DE8��b���-���V�R���ǮM����ű�̪O��� q���C�c��2{�� ksc�	��!�sAh��W"��>�:\u~ �;��f�P�j��ږ��b5�}�~vf0�K�k	�[�R��p]A&��TE�ً��kҷ+�~5���ys5�<gi*q+�(�bF_E���g�,E},msel�&.�%1�c�*�=OEƇ�%[H齄�Zc��j��x�'�enr��*��Q�ǰ�=��C���
���P�#��	����C4]Zz���)7�(j��`$*��������H���'&]�9���x�S��,�g/@�N!TiЇ�2��YM��YM�F��c��t���`�Ҷ��_��ȇT��<���~�k�TԠ:�BϚű:��IF�o�x�n����v4S�t_ja��7�;��'ӂ�I�A���JT&�Tk�z�-����Őބ�f��{�!��22��%,��q��)�'j�w����ێ�\\��+&��s�+�S?X�����f}d�L^_���`"���ә�Q.����Q�>
�t-�a��9�����S��ab[���i� x�7ߛ�4����Dt�\7��_e�nA ������7�{w)�Jܳ�:��u���7���77�Զ�nJ� ���k��*����|kX!P�P٬��e5�3(k�o�-z�Ǖ5�R��:�����]���Mf��{���H�3�ЫE������ZT�n�oe�>K�]��o�Y��drxa��� ��������2�M*o�u���8�̀c[�.Ͽ��?��Lc���8��疚��D�O�!R�=��i��ݯ�n'o\
��:{�\$*�7s��#A��û@�b�6�J{m5�m]Key
׈S_��� �o�']<�mAi���9[����X�r���NaI�6񡺒4�_j�q����q�����Oցk�'֖@� �m�'��t?����N8��z�������Tjef?��
EIG�8n}z���k�%�Y��(�d�c�D���5O�L'�2�e������,���+� �0�gT�m6x�c�i�+�g'듴�&o�SyY�o��a�6o#�T6�e,�y�2O�-���Y�y�VM`-��?��RJ>�8wJ�����8įv�/ C�6<r�gn�)���㇫T����-�"q�o��G"{G���i�����|�0{^�$T��� �1�V�RN*�60Q[k}�&�r��y�x�b�:{�N?�gA��{�1��^L�"h�45�l\G�}W���Y.g��g���R`�����z�$� ����gn1�6l"�4�`�hV{�>HB^����ޕԿ�8ɭ6)%P�,b�f��ЋH9�~Uf1�H��ڏ���r��4%Pl? a��歹=?9N��X�3f۹Q�O<�� �N��g��[j�.�1���{�K=A'+��L������C�i
I���W$��D\�x|5���y�+*�A]F��f#b�����n�2�(�x�ؓy���,�/W���5,�>��"K���O*���`��ri�z�Z8"�:�8Y��^>CMD����� �A�qn�������K킄�-�l�{��_<�[��OZvP&Z:�B�fK/�<��O�ek?�J~@c�9p�c&���d�0��J��&m�n��N�uU��_�r!������~� �:��+�z��j����w˨.�'4E�����W2���$Pʕ�9��2f#���R��T~PVs���R��aǾ���97d�����G&�^��
5 F%���ڜ�imD�J<HF�<v8�!�0pر�\x;��!�iP����F.,80٠y:��[���[�E�xN�U>�?~<�C#���u_/�&#jX��r�NY�Q&�ͦ��k
GpH��SH�R��~e5��xR�ͳ�b[�D��sV�U��rΗG�?�y�s*=�M�1DrE��ݯ5��{�JK���%�l�	���(,�+�����(%��9�d�&<2��~J%n,�+	�`/�Mf���'�2yJ��gz� �����O)�4�B=T��M~�y�Ӓ0����"�}�G�5��S!J}�2����n�y��^��鷗�3m�7��Χ5}����,��?�������E���P<����d��vN�L�?m�0	+�vCǍ��5Abq�^�����E���E�NK��m{�\"%!���5��8�j�Y|D�F�[�N�!�E1jJ}lGm���:�4�й��@�p-S�����K���T�c��8�.S����2Нb>�h�mX(5��c1\�;�w�+��:�O�u��Ԍ��}ևxݲg\"�l����r���q���kO."r��V�sѻ5a�mT@YS����j��j�6o:���џCGp���@�M�����9;���+l���y�7<n�Kx�o����8��3\��p|C���k`�n#N���y3zc�k�9�!
���i+T�	���R�x,�P�����}�&D��A�|{s����B�\H�5�2qm����N{�E�����M钠�V@�8��w=���qm���Sx)��{�мW<Z���5����5n&V[�@RI'�5̨���Gl���˳�a�v��Jz�C4���.'��x�ˡ#+��9�j6�r6n�סM���k`x�����.�����5�>�y�, S��������T���O*O�(N(y�K%�hO,a�Q2�O���5�E�N�ѥI��87Z�6�NtWݙ�٧C0�6C���#3	z�X�^&ڤ@8�:Ȟ:>�e�&;o����UvEL�Gsm��6�ʜޏ���Sᔧ ��D���T���������W6�8�W�P��/
�=�W�����K�h���,k�wZ���3��"Iaq�w�g�>'��ϩx��f��Bq�x�P톪a�� �\���l����`q��_:�	o
Jr����բ�0��;d��H9yîFW�7�z%{�wt4{�1�o��v�Iv�	(�� y�	7f_�`�=�-���s��6cIld;����"�e�˟Gq�!%2�����jf�N����29��3̙$K���!��`�I�/�@�ki�����S��7��	~u0�7�0��y�D�y�~ؘ/T7*�s�b��>e��Uu��w�%��f�m�E��髇<��E��_��T���RHrg`{�j,�C����z�V�ZL���F_����~FZqe��C���!b�33c�O�M&נ�\�-����ec���Sp-�V0D�W8����Q�}�(vfW@�)���x��ͽY���瘤i�}Z>ǃ	�w����!�D"C�	�z&S����.5�ȱ,pa�7h�\M������4$A��=���l���I
0l�������򗺫X�հE:�`�a���R�M�����K�墻���UL�Y���� �Z��88�k>!�z�\����� �ѡ���ߙvx��R�02�e�39{��Cֶ�@�� ����'�V֓<����3���^Nu�5v�P����M��	/Y@Vސ�'jH�_�En�3c�Մ��C�d1�`8O���ۄ�%QLr����s�v9Qkl{�O���$������[�F#�|T�)��`�""�]�#�xD�em���Epp�J���0��h��Z?|� 4[���j���c���fÄ�:���&����UNxޣğ
�k���泠�8G��5����k��Z��Hk9����u]��؋��?��j��)��!�1�QI����������v��ί�V�)�̋��=�H�g���*�A��L�߁8�u [i�;}�4��A��8��g�7��ĸH<�0 �2�$g��ҩ����y4�]��E�i�L>��P&�+���,H�����̍�|���Ʊ����[�l�첮��f�<�W�N���e�RM/�d#�� Kܞ�)�Y1㋋��������f��̵��_�i�+%����,x�G1�2>���i~:�H���7�Q,� �"�%nwӠ�$[��H����7tEv���iÚżЙXM��G[����F��JTgz�d�@�!�rvt�Xޚ�2��|�i��=��8�~F=u���	U���W�s�y>���������(���B�"�K�Ij&��@�ӹx�睊�[���8��B��U9�6��4^���O���$&��O�dp������p ��堳��tO�2�?Í��XgH'��Jy�Wՠ�eX�Ș�{�ވp�D��Q<1J�G<Nm��6��
)�Ԋ�\��z�����;@@B�)��ī���Y�r��>{j���~�A|���x7����}N���=������#��	�0�":���Q�������0�o�J���Z Zhm�����钡%�F�����1Y�"}�*��6T��uT�[�3/b=t�jP����
%����=���|p\ �{���|	zs����� ��C+X�K.��0Aє^�-v�^EO�s*�\�)�ˍ!�@w�z3GQd:h]�'�t����^��q"�:���36���$����5o��Q&�Jh*�Dz�+�U�i��֗���vt��F����y�Q�?q-Ɇ)^@�"�\�J�Ȝ��ef����V���Kx̀�}eV��ȧ�O�%�n���_$Yo�i�H^�Q��s���k�h�Ÿ�}B���9����Yd��u;��2��3h�y{:�u 8�����S�D�"�*�YQn@I��G��E���VffA�ꦦw��]�Ҧ����+���Ӻݿ2�F��Z���� �20���I�B�k�<Iٽ�����A��n�=A	m<���`#�]�LՁ}���O�A>/q)����1�m@�LCz��@,D�OD��)-�e�a��{��<���`�F�d�Mr�m�̧��MT��������ho���Y��dm�5��RS3�>Va�R�����hCٱ�0��&�9ͽb�;��BD:���<m�z�g$&,��Y�^��
;x��e�<�k�1��#�7��uT�����N|ef����W#���/7�	�a�9�_pA{9��	�-yzϷ$� �R�O{.��mӟb��I�w��sC�������V0X2o�����A�����&^��U��
�o��&>{�g�b������'ĸrƌ��	�Գ��
���t2��{���c� �3�4)Y������)բ���X���BQl�� ���:ׄ,�����zۋZT�Se`�2��� ���d��J��{^c��7O�����Q�qۨg]�6�y"?a/X ��6��&d��I@<@e�t��vl�ճ��H0?+~�g�0t���V�U➥d���d¾�۰V�q{U�޴mȷ�䛅�A�H;aN�n�n��C�;���j���8�;���a$RYW�M�v�惙��FMsm%X�r���;��uaQ��[q�dK�In�t �#le.&̀���Ű���j��������u���@�j���4H&�%|sg�m�O]�)J;��M8ڮ�6�!�(��6�wa������=��$��?�T��2%�%���<�Μj.�������M6��� �y�neDu�h\�S�R�Dy~� k%�a喱koדA������ʸ�����'�-�D��*<�Zy�ڵ�9C:_O,ZȬ�W�n͵��aQ+��/{��&|{&�E��[��<�Tq�_�η�Y#V��[��P��� "8����l���}U�K��K5�ta㱵�$��۹O��"�hY�l��R.�g��zez+e�a�{�C,# ���#h�-ov�BX���ӥ���b~�a�Z��8�$jGK$TF���[7O��C �4�������_Up������1.-q�ϽdyFS�Ǆ'C>+R53�VKxeo\}#�Mb��ɿ�{k���;+p�����/n��A���)�aO��3�#�R�7�a F�D�K��	fX��뒧۸A�%�'Q��iT���>��к�>I���Ґv�<E���&62z��UI�v�>��->�%6އ�~�%c���ȸP�Ʉ����RqC�2�QS�dPc#��'o�����S�%�T诲`0v�1�蝎�v�1�\��`����z���dм�ꅊզ\޿թ�|���>욨���y���Vd�d!�� S pδ��2v�td�V�������l ��@+|�#�g��L��3�����u×�(����'q�K�=����{���ʢ@�L
#] K?K�d�n�;�����
��C���N�9X��&qCz㣝�E��f������\�Q��4kf���~�����Q�a>�[��h��^Yߞ_�(����~�j���I�R�����;4���y.o��:����	�3���� ���p���]w�����F�䮘P����P@`&L����1���o(>?#?U�U�\�K�c{m�U�π}=�?�b�mW@�ک�H���/���}�>g�s����]f�q����Z#�H�7/��=���	���M�.�o[n�Go@ɴ��s��(`8�F���4�?��̉���h�o6�K�3���1����"�E���n.���f����E����:?�9,��F��>�tmE���YU�����l��0��@�����n�N{�bGE�Ǻ"!�� �X��s����w�@j�J��W��������p���4zZݥ��Y�2Y���.bp<u�{��8�7�Yƙ�c{�H�"�D�"�,� C6RT u!�[a��FD�V��m 9��p�.��-�#�`�Νi�7Y��
��O���b�YR�����٦�fY5C���[��VS��ͅ�q�V�M��'YJ�	��w[q~��޹iD�������KA�� 5���b��y�T9OT�ȰV,��^��V9_���}*(ˆ}[uqݐ^>|t�`S��6���C���r,z���`�R�<���p'�0��3MHc+ 	��Ԯ���G�EA�j'�s���tڈ"��f�H/E%�,��e���	ZY�3&6s���p�P�W�5\��b:bi�C��w�[(_x}8���䲕A̒�4�K�����a-���7s-GK%�~��b^�s�2.���el��oư��\��p4�R�$5�m_�Z�V�eZ�+�r/W]M͝6�H���a �@��$��!��8�C�ꨓŞ��߿biFA�J�z�|HU�j���7+*C(��"��;:w��Ԗ��>p�W���X.
ģnOT>���ך$�7�>�n��NB@����a�)_1����
�P�jUX8!V���(`�����Ц��R�� T�A�'i'��O�_�����6��#�^G&���>����!�ÃTu�C�9�c(�1F�'���Uy1�b�a�����u�4��~N��&q��~}��,�j=�+�0�D��I�Rl�$�`�91)\���kv�ֵ����������(��7�e�L=��Q� �ΐe���Qo�	A�[�R�'�������U��b؁�sE����������L�7ז�ݞ����&���4��IT-������Z�� U�gQ�ȸ$HY����'���3jf���&��pK��9M�s�`��	!O�L���"fJ[��_3�-�f~�Z���t�噐��zh���c�/��
Z�\$f�\L�)�7��/�����{��;���v��{�$�?P�$J-τ���9*��ٍ_$�TTFŮ6�u��=��VttĜ^܄K=	���]���'H�/£���p�sl�����ya�\oer�`��w4���>��8����3|�ɾ��<:�O,չ�}x��x�y�g��2�+��<��K���L:yY�����K������S�)CFEQ�ʿ��na݊�ǉ� C�=���5�|$(�����qfAM`�F�
ȵ��O�n}�I�/s�v\"3�M�-�X��v65y|`-�����s�pEE�є�O�q�̀��L�D�"���v���sO�1�m"�R`�Z���	z��.���U;Z�
���{XX�N�^ ��{��Un�U�|H������*9�fe
U33m��VS���i/&B]�HjǤ����d�^���:�=b�*��Y�K��-�I�=>r
��_8��������댾�rq_E-��2Q�KQ(��9M���"����Z����� į��nU���g�̒�%;���Et�S��d�돛�X�-��i��ɜ!gxE�|z^Ʉ��8���t�@��M���Ll���)�d�`�㰉;�Q� LEQ�)J	�����4���&@�!�w����v�v�������Q��K�]i+�$����Z��wa��|gL��ZO�o��F>r�P�@�s�W:E!_���/�>O�O�b-���N��y�<<Y���]���S����4t�a�/�TG�Iz��P�%�vJ°@x�g�����*����UnXq����s���8��^{$�M��IV1䬡?d���@��.a���nɬ�O�]�\S$�mH�/gE9��4��`'��>�?*vn �y�_���,wj㥃����t}���%�c�s\�����'D�z<:a.�ɭ�C��`�+���,_InKq��e��2��*��k���?�L˰��7�8��m�Q�꼫�`i������a>�	F��3C�~�?��2�`��[M��1�k��hI�#|5��[!m�~G4O�9�@�����h�����B��=̏����2���ٙ2kj��K�M¥���u3���m��:!3������Źv�"��p� D�rA��n
a�C�7��7�׀��p����^j�\ۍ
��(t���S��fױR��BH�g׹�r9��&����?L�fQ�0��J��j����������@�h�i͟��g7]�L�T`��	�i��2E/��kE��m�fwu�'�E���2(�lr�����b�l�>[[�F�����BG�F-�U��n�y���"�����4~��a #|���j�󱜢�#��������zi���DΖx�؝"�?��p�D���;���&�k��LG�F���"_�# ��!��O�i8&~��;J���ƍ:�b!:@1hff߭���0U��p9}֩�̠���:)Ci��$�U{���a5�3��cJ|��X>'b$�p��l�4�)}O�ڼ�z�	]�1R�ǌ]��y	�t�hx�՝�
����N�� 9%8Z�8��u3���Z^�m�L,mH��r袼��4�br�(~��rp,9�F�N�'�M��_���:�\8V����e��\Y(<�(1�M#Rz׸i�q�!�ȓ�e'��h�-� 0o��<rN��?p�8�z�	���]u�6Ϋ��>�t؊p�f����ʬ�8Uu�3;�X��?�{-�dI��C������ ��J�cUHHܩ��ik۲91`|O���O�lb}Ϝ�H��`�5����"hk����]��sge�t��V�nrd����,&�̿�y;;����f��tf�,�y�[�N��71���<�-�@�O�I@�cGn(4e�qJxñϢ/��ӥq�O���J��7�W�
mƇ63;�[6��tmF^��{��7?�ڻw�z�݄xV�F��j���Q��È�})ۏ�|�+X��Ʉ��t�Åy\��B0���=�h�	;C�IW�ۆ��f�-ӹ�9���zK�}�̖��g��,r���z��ֽ�!�7<�]����I��zƣ�"]���������㩇\��ϿQ۶��n�bщ֑����>-�_잳���}|C������n�@۾/vdJ>5kp���"���|�J}�f�{ߜ��4���а�I�m��Z�"K�&��{h�x9��B�P���y�3����S�Y�"yw6��.jE��cfX��+w��Q$�߲+[�tS�r�{ǁ�5��Y�kkz� �I�`�,�H��!#!��l� J7)��Jlσi���X������`�+2��菜�"�����8�Nօ�,G'oM��u��-�z`�aq�x�(��^��g�k��;&�ܳ�5x�,�.����hR.�^���Fͻ���	'|���I��j���G^��R���Ɣ�9�!Z�w���7��/Fq�>�v���ӧ!R���G�N�c-�X�tVE�����W=J�:����i܊�$$��WQ�ı�#Y�����f�B;5�5Hk�m��2J� �8w&����}��@�ԛ*lm��.���o���,���t�B�rZ~�?F�,��x�o�du�,��>���]�P��3�\��$��㶅�Fڬ����
�`��5���`���o��+����_��+�e,T�촘m��x%��c��~���}Nꂪ����-�����3���7O��vf�MY�^�Ǆ�́�G#�/��k�|}����A�l�Y	N�aᇭ�Q ���s7�n�\�(��MTEƹ=ц�1c!�o�Hu{��o�� hOc.���1]2��(Cr��v�P��7��|��ϫD rvYq�9����p�4!�|�g;L�H�+����b��r'Ә���H0#��8Gl1s�ۏ�kc�J_r��I�A��|��e�����ڝi���rcRr���Sk8��fn6:�Q�	Ȕ�&뫥+�[ğpޘ�QB����j�a}�� K�w30�8��(�U�9���fha	Hr��.#��;:H��Rp�)�����(]��B�*[6�9�ƫ����M���[X�W��ܕ���j�1�ԭ�9���<����^��]�ID�W�+�zf���]�+K��:QK�׫�eC�c'��'cp���ܹi�0����5[j�9�4}Ư���S �n[H(n��l��Xps�ѷc`�a7=��^���֜oߚ�b��t�U�I��i�Y��Vp�/�SZ<�������hc"�_���x�&���{�S�U+�V��G��v��u������to�8��mڌ�$�i�ʶ�_Y�*x��C�,��97FF7t��@��c��&6��Z����Ϝ����G;�ݳ?[￮�Pi�y�V�}������W�[ήu�s��\�V�M��������O�4~����.0��d�����z��f�{*t���k��'\;�3�^�*�^z���k�#���M�r��.��3#����o?�gdjx�ND��������a��'�_����	ۇ�'�R�xP��bDf�~�n�R�58n�N�֧yLZ �r�������1IV�!P���i�����5(��6�!_j͎fr�/MU_L&�xr��,Ę��j�Et�LU�G��*��O�ЙJ?zq+vOL����O�>p(�LX���9���NK�v8Φ�>o����9��VI�!Hĳ�����^�>*�]p�5���VVJN1��8&���m��RUP��k?{����^�Y��.u;�n廩	�6�vn�z(\�J,UR��i�6D>h:��=��i���H���G���b�f�tR(��_u�;�	�1��R�uZ%�#����M6AQ>�����2#�~��vT�y2�8�&�C�.�:��)<��}~赹��$��X{��������
���4�j����l}�?�p7��l[=��M@��'�Ƞ���6,���sx��~iD
���~I�����?=������>�r$ܳ��OX8�����,}t�������V�� �� PK   �n~X����}  �}  /   images/e0206f85-8494-42b8-8b98-142c319be1e7.png @@���PNG

   IHDR  Y   p   �&�   gAMA  ���a   	pHYs  �  �(J�  }uIDATx���eey���]N?3��� Ì" `�c/�c���h�o0&۽��&�{cb�o4�X�l��F��Ҥ��3g���������k�g�}�t&<���W{��}�[KYD|m�Z�$��j���N���9W�T����{��E�)�lb������|�́z��Z��k�J�7�t�|wn�A���6Y�����fz��G���Ӈ��b����'��u�N^�������?�
��u[�v�5�M����F���V�~�-�6�p�@?411a������n{gA����x�:8~�i�={������ƻ)C,�W'��ʕ+}������ի��O�+V��8�'��ܹ��nڴ����н�w|���������~�_O�1���C�K�Ɔ��|��pr7Z d/����⋽b ���h��633�����U�C�s&¯�ʯ�߸�����|�e�y] �3�<���������$c���3�X�L۷o�ݻw�޽{��Z�h7���O�rjъ��h���s�mM����j��������=��2q�����o�/|�����l�3E]���?��;�<������������g/zы�I~�0��Hs�yr����&''��,/�wr���b��]�����&�V ��k< ��dr���������-V����������mo{�����g<�644��i� ׬Yc���=�yO��2��w�9"]+�T�M;}�3��7��~�$\ó�� )%^�T^ ��������|�����1�����?������>��O{������^���u�]g###���<�n��V�~�D ���z�=��O������W�ڎ;���Ї>d�V��w�� �a#�6��GZt�w7.r��xE��Lr� �����p��1��`�<��ϵO}�S.N�:΄���z��^n�xǟؓ��� da��_��Yy�d���Ȟ��g�_��_x[ x��k���?����u/��{�ӟ��nړ�<�Ї�_��_�'?�I�]��9������g���E��pM�q"5�to�v�rN�v+}�9���)?�X� M=OD���%�2��^�Md���gf�>ƹ�:|��o�����lDR�J�9���@��PE�Ȁg�r�T4�˖�^��E����ޓ#Có�3))��Ĕ�4Z�h�mrj�v���;v�`��.`��5:�/���I�}�z�?q��N(���m����խ�v�R��gڂ�r�w��7�쓗���:h3�z�1��8ޣ�ʜ:����)�~uЮ� ���^����U�axW�R�Р����1�w�vZ�v>����CEb(�t�'�t��[�����w�i7�x���D_I�twW��,h��p \D�h@�k�q���%��n�B��G�Ӵf� �վ�y����j�
*��e�Z��E �|��B����X1b�������3�*�7�s�_�	ў�׻��fj�X���a [�*�Q��8�9�O��|�.0��9��E\D��q��b�H!���I8~��� ۉK�aw�v욵����V�\aS�gXP�����<�*�@֏��G ��jq��I	�ޫ�cuW�=s�>н��Xړ��9�y��n`&���6�����C*��<��NT�,�|d�@�H-L7�
�&�V|����1�P� ���d��y�ѱ-[�X_�Z�l�0\�9��������Ƙ|5m�s�����k��M��1�m�28�a� ��uOફ5 7	�lj������;i�[�z����=/g �]��|H+?���12�<2Щ/�1���礃/��Ջ�u�HN2ѳk��FL������/�5�]a�������}H({=\�Y�Kz�]������٘����4�?�~�e�m3��V�j���w�q�;,�M��X���.h/��J�s�\,e4��+�գ�o��0c����L�G�v�� ,��/�+s�YC��l&1`��������*���x��AJ����t��?x��v���#������Un�Ȫ�Y��\5��VxQ�
*��W��rtd�>��?�`�AH��
��O}�����u;�����^wx\+����خ;��&@��L��F;�u�����7Xc&�ch��պ}����2�Q=X�qN(voC��=�~���u���l��ڳ�K�S��<D�Q)��ϱK��Y`J;Q�Xo�w��+�r>�֯_oOx�"��ޅw����	��)���m�7���XX�BY;��7�2�G��pEa,TB߰@6��ljl��Txw%p�I����nb,��,$�l.���C3��M�#q|,��W�
�9���\'�f��\�$�2�Ɯ�b +�$$@�x	�֡��
�e�oR?>�y�󹁝�^=����t���E#�:~(ݳ�4��i��ux�L#�u{�Sg��>>aź�����vML��}����TҶ�^1l�z�S�� ��9��|��g\���Īu�}�sҶ��G��?9�k��x+��1�����_��pe��8'�vV��:X� ��<�)����ۿ��9�\*�i�Įt1�j��3c�_���{b�{��]����]q�~�����H�Z�����>e���6=v��o�[��XE� ;���V��	 ��n���	����N��u��+Sa�>���_[i��΄����UO}$mY?)Д?x��\�q����՘@��8��Z\��x!_��
3ó��Gڃ��b̰�nܸ���1�^z�.������\m06�ˎ&r��� ����������:P�1���W�ؖ[o"zӁ]���۵�N���BZ֞������׾��@E�0�r|�.bbZX��@P�f&�_\f�V#�O �ڠ�8��v�a����;�=�����}�^�����Cl:��c}���T*{q,���KO[�eД���dx㯀U�|0�A�`r�%+.�Ƥ��@�����i�Y��bӁ�,�S�� ��x����X��քu�v�^"k���Pϛ�^Rͮ������g�.T��ﴈrs[\�8_�b�uه\���2������/T���r�s�ٽ���f^��b�=�Q���.��M�,E�����\��2�8�XM9�A�kXc��P��(�o�8�1Y;&M���f����LO��7]�����-L�0h�Y�"W�`�9 h;��3㻬ڜ�_���0tb�U���l�U�ٛ��f�C����n�C$Ql��Z1XjR��|� ��$P+���5�{ ;&%ܭD;��@D��K,<�x������-~V��O�N�H�?i�hU�������f�b<~}�|�� �m%�T=]�G���$	@m�� F���P����W���h��7�v�W���2� U�S��9��''�Cy,~R:w�}��� +�@:�He���?\ě+94��&����L��A4
�H-�g�dk3
]-��پz�j��L��S�}�uҁ�<�K�yG�����
  ����]��;����f��#=8�e5�~�9M��bs;|g�K|�39���*����w0����͢�r�^Y�¢�I�Е�@R�0xF�k'[���#�F��
�F{�_;iXt;��p$�Y�� �~�b^�
G�)X���� ����,h
6����!��b�i��.E]�;Y���{���~�q�#�.W9�^�(wwr�e%��u}G���L�]ہ�&m=p)�o5·���T@�D!�H�����d�CAY:U��rn��	I�iv4]��l�
�f�	����pAq�g}Wv��"���b��g�&�;*�5Y�[|M�����{E'�j- $҄�Nkxu����l"p��J����J5�YNh�0*���=��2��H�e*�إ.`�`D@c�c /� �b`��<ci��g�Bed�m*`�u��g.�h#G�4����#��R�.���j��ИC/��x��N5L¦3�%n=��c!3�e�ũvE��39����}��X�	H����5�;���p�.e��\_�KIY����.�sg�wx_"i�T"g}��p��w�捰�ͤ�kY]_	׊�Q��N�pp�
�b%pV��a�m��j���7��G2��U:s���ۨ /�Q��h�f�N��/����r��cn���cgǎn��֬9�0,�D��G�y�f;��A�q�{�7��~��Y��h�w��,�=ܽ*uSE�\�3}.��m'�ln'a�%+��K�01�IpA�/��t,L���Ybb��׀9&i�2.j�3}�k�)e��^LӺΠLe�=�&����V~��� @fP����(ڏ�	 kᅤ���Ё�R����U�.U�_�ծ�Lk��L��¦Z�V�ΰ�H&��˕���]����WY��� �j����6	@�d>�tm�tͫ28�9�4^�lU�}1.��D���s����Xz�:A6I�Դ������w�~�||]{�v�9��bhNM�8����"���aG9:<����dT�8�+��bVTՑE���i�B�6:u��kL�"����	���g}�A|���VknUNj�a�N�h�h���t�ډ[���a]�Z˕���F8�n-
siu^��^$]#��rIj��{�����h �@@��� �Xw��������H[N�$άW���+C�����N��>���T�_���n؆�狮���)L���\ak֟� >���H���I5�a��^2t��#T����N�i��X ��O�п�\��P
8�6)�Ȗ�i"��_�җ��#e@1�)��C�C9�N���x�5cG9��񅈁�0Y��l�K� �@� �l+p�ͤߚ4;ؕ�l �Z����W�e�n�m����v��3M�E�V���L@�F��>h�� �\S�6�A���(�|��Yy����F'����� v�M*^�ԊQ<�c���I�#��Y�m &%�^�tuʛ �#/�2��
4Ir+ˤ�1
�%�@�>lë��k6�{��Р�w�񻳶�X�����P�����kl��4,�� ԣv���m��v%���=2I��rϒt!OڑvSv=~C��3�IB�z�Ֆ3�AK�hU�m����� ڻ0̉�|��ַ<��јo�A��`գ17m�d|�==\Y��|��b����|��[����9Оr��`3#��R�P���m��f`[�W��k�%��fbh��ڥ�_�n`yO��n�o�*�!;���u: sÓ��<&L��Uw$D���1؟�ԧz:=��,�d�Z.Iw^��k�џ�Sj&�\� \���-\��Y�)�,㈲���x�Sf��2e�r��,5۱s�}�㟲ϯ��5�&��J��J#7D���?������_`6�%_���o}��v�����q��\,��?Ł�h�/�RU_���/�	d�,Ʊz	�9��;��Z���7��^���{�9�P.T����쳟��/
�:����Q�_w�mݼ��=�\��W�:���b��C�ɨ�4���G��^q�eC��7{�{��k2],�8ӝ�m�1� In�]9b{��?�d�)�F8�GV�M��@vڹox���ժ}�_i�ԟw��d#�;��gq�3۹{�V��9�J�-;�dx`З���Ջ�D�6�@"�#�$Nj�XJ_� W_@q�=_���A�:��P��/@@�x����x��69>���X�|�ߴvcƃM|�U�X��;���@���O~��_�=A���6i`�I��3�)�Xo�j�F|fVW>�j�*;�ږ��TQ]�wY���m1��/�1�.��J��_�Wr2?��w�	��[n����_����1�h���0����۶m��s�(%���0 ?;:�T~�Z�>��_$a	��9PW�D���}-S���;�/x��>��
��0�v����83^�9І�������ăjy�FGW�W��t�#lb|�	i�V_�M��_��LNx�ku۲}��֫^cY�IN�!&H��r"��X��ka��a�ᐌ �\�8^�W�ƀ%Rs���-��P�C94^x~/N����"��(�[c�|ǡ�C�t��I�s=w� z���� ��z���Z3�Oq�!� @��J&R	P*K+���uYTTѾ��Oٔ����W_�X�|)��Ƭ$�N��ʧ\Cg�z|~�t� ��>�4�,�y�C����o�l��E�F��~/[����}�;G��p5W^ye@����̌5�˚�<�I3~�&ؚ2�\�jxgzB�=�*e����,Z+�`0�>I��ڲ�'*�;<:d;�NNMg*��o��xh��ǥE�8b����/�&�H�/0��i��sqK����Y��L~��Bf��N<_��%抓�3V鲗�<Z,X�k$;�;��WH���m�3�=�}.�dYŦf�{ZHcᙍ�5B����8�t�uٌI1�k|G7�~W.h��+�&�/��
����_.�R*~�0q��r,���I;��V#�'��́�b�n?��O�\�IB�S��Qn��e�D�x�4�-Y ��:�u���������p�&�R/N���Intr���p�2G�
��DEDL7�t2�V;�lwr ��T&�w%E[�&��^϶5�j���hF��̸m %;g �(qN��'�{\�b�x?0M9���_��ͻ�����-�j�1"��{6n��yw��."#�a��BP&���< ,�㡯��\g�������Ef.�1��)��{�}g�ߴ�_-\K�C��?���fm�Ze��u�i\��2ȱ@�p)�E�I2Ubq����c�������� mL��8�*$;E���]�;�`j��|��tӍ���_b�����Yd�J�*�/۲��E�2���x:���\^�җ�s��G\+�^�f�F��A�ج�<�я~�����g��		s�c����K»�<��b�5�3�$���	1����j] )��=����E��;e��p
㮣��7����p}�!D��v+��x�g�_�'Zm�����b�q�8���{�����~�|�C��20�:�B"ρj�;�m�d��aa�ܤqTn۲5�Ԋkj������UN�wQ�'���՘>��Wj$��5�#�������?�3���Y�<��pj+Mt��������?���^���~���(L"�����v�eW؞�����뿶����jX�[�����v��?�A��;��-���@����H����,�d�g���R�t� �$ �A�Tp�ާ����F,�
�?�|�%_���#����I�����l{�<1��Z��ٲY�"��-�؄kI��%A O33P�dLN��r!�t�{bk�l�殫�鍿��)/�3��-������w�����׿�N;� F���3Р������'�o<�]�`�)"��L���=ا��	dRV�{��_�;���ԁ:�������Z��o�ۄ�k��d����b=\ٸ��"=���h�v!lz�ĥ�XT�O�UA�d"q��->٤����_��_����)�mu2������;>����ź���'\������3@�xJ�a� �4=z,c��;[��z.���K��qw�kDj/y�h2�� 	�݋3�#�bq���bU��Jt7c��~��H��9+��ݻ� ��� �-����C�}�M7�g�^���(�Jᬳ�r����~��_���
�=�&#��I�U�0�y��{8�l��Q��׿j����f;
ei������é�*�M}��Z��q�vpї�h߹��������n�$�[����pHB�!��I?��߻��r&�1J"������0$�Wje�*�K%���
G���� �H�ŲN���p��ǻs�N�H�|���c�c?N��~lm��Q�}��Mq�<���{�ě����5�$�@�.�m��Y,�k���ғ����qՉ��1��nŹ.ĩ�@����'���@Ώ�I�u���������c�,BY-n�NdB �p�tp�hw��dp*8�+���Q3 �sLz#8e������F�J�:rN�("1�w�_����n/+j�һ�h�_�(��T�t���]nM����c��db�ws%q��ń�'�"�bY�9����}�X�O��f|'�����$��/�
�е"����>�����
�w�]���Au���i-��;�\���ߏ>r	m��KSy�\j�k��x�cڐ�ߺu�=��Ϟ�K�$/����y)t�g���� y����a�)60:l��]��ozK6�;I�b���(Y|�ϱ��R�)ZG�ٵ���݀��7�5��V!���]��T�EO ��u'M�MJ����=�O�g�կ~�;W��EU����o?�w�����m��I�������}����&������Z�ge�P�z��%Nm�g-RjGE�R��.O���b�e- �N�)��Bnw�_���RH\�^eKr�T��k*��w�>� ��|b�͖�h-���3�V�O�O��fd�:6�v�<o�mZ-��q���#�b#.6���'����p�ُ�5b�r9�J���x	�y|��_.�����a2� L0�G����]w�� �x�qq<
�C�';�s�i���,ʟ��d�e����{�R�z". &�ܾYc����^�1�c!W�p�k��r�J)U`#�;4�4�� ���c/H}��ye�,F�\�1�/F^�����M�ھ�M�@[��b$�1���Y�.c�1�!��/|aΕ���ݷ�qK^ <�,�`�C�}�[��#��#(����!�HVi,�j�
�ܷ0�UA�'��dt�����4���0D�X'+@`	N���<��H���?��?�A�j{r��P�CdsŠY���7-���� ���?��.���Κ�ϕ�7׻{-���;��N� �U�z���"�o9��qy1��=�W9	���6C7'B��g{-��\.`�o%�-c!ڗ:.���%�V1Z�ō�M�	1�q���ln�����ꝃI :�^TI��<�>����`tx�З+��l�)s�,�1���Y9	M��� �3`��T��+�2�A�����g��Ā���`ƀ�p�X����A]�M� �#��'S���8$v�:wz�P(�;Uĭ�9�2�L@I)�<!-Lz� V��+DV�GV��-n9���n�>C�X1��z¢:��@�W毲k��b-�w�w���%��iwk�K�Y�>mE���\�|T�>+�/���͆�V���F��tڶ��f����%x�Sj�y���l�����[��d3��ڵ�i%ɘ�i�yR����~g�<��1p��g{}��1b�e5��w�ѽ;���.���}�ۣ����=E�z�3�]��$G@����?��x`�`[k��1ɐ#�n���ҥr���Ew��hƠ��V���ZC�|6 h�����bVe�Er~�G����O�J��{�V�u�0"Dm��'�-��6xi����h(0�-�R3�H�b��#�v�?nW�!���3��Tʆ�ʘ����F|�_l�����v���������5��7����w�����>l�������g�#�����Vz.��7ߔh!cZ��`!�����>����"����h��1�L��6X�Y%�����l���ju�����k���l��z��_�M����:�tn���N4۴r�m����V�����C�pjY��u�N�X����s��|1�ߩ #�(�l%֕�����Փ��R�D�܀�(d~з�2vHܧ��I��2wp�y^�V�� u�L{(��8%�^5\߮tˡ��k�'��s��ґ��Ln���T���$N���Ї��DT�/��e�� b#D��^�"��2i�DZ�K�
��J@|ߟ�$˥^ 9����\�������X�pũ(����eD���� )�9�{�=TN�(� ����xJͳ/a�g���{zIj�b!p!:�*p�|�h>�Q�{�Z��]:t��8�_��XLg����E���-�.e���XW�8�>PN؅��ُ+��Lڎ�.�mw]a��������b���g���4���mV���J�P�8���7���0�UR�B���h�e�]z�5gP��XN�8��2h{������ɛm�kent��x"����}���<!�{/�mv�WىǞi�#+-���m���p�Lf����k��?��μn���A��M��y�U?�Mg�j�2M�v�{7ۺ����e�����r}XA���[�>�?$<40�|�K�QY#NV�����������Nd������ØR�q}  �DDY��LW]u���=�iO�{���>ix�c�+�\ ��J�r'ɾR�7�yfNP|!c�;�� � �8Q�6ѓD���;�r"p���Q�O���B�LL$r�|q� q�j@�Y�!�L,��|�+�lx5��\���.r�-�e�� ���W��@:;�L^��U�������']�M� ��o�7��	��,Fd����js��[1cC�Uۺs�5�Tl��Uv߳�U��>IMq��,\\�O֒�V����,����b��7�L]��薇+g��v?���p: m� �a�OWX����g�9e�S�|�PCC�C�t��Ɩ�b��~ӈ��������Ԧ��n��:;�O�dϕvݏ.���'��Y�Z�o�/~�C[������������)����f6������6����>̦�ή��r[w�1�?\{�]}ǭ��������?���w���J�|CUͳ���A1�3����-	�{:.�����ˠE70ro�v�k�ѱ0�^ܘp����X�*v�I�����t{׻�c��h�:W/��.���ќ�zJ�=�A�0	���� ` k.rL��_���@BmCc� ]nl�C1G�ꉈ:�V����yu�|�D��D�l��(ϖ8M�چz�/��x��N�^�g v̕���˴��牉rc%"�BYL��X������&d1r��� �ɸ��|��~�����+�\G��� �ߎ>�spm�g8��;��۾1i��q<ie�$ڐ����,��o�����]y��A"�@g�M�]m�{N�k[�jp��]9f�3Y��*�p��K~i�9�j�%fv͓�o�=��;7�u����8=p����&~a�\Ӷ3�촾����{��t�����_ص?�Y ݍ֜Nm$����r[{bx��vk��n���)��Ǫ�;l��?��M��Sv܊������m�����B�����aλ�/e�I'"���B����&��ie����n:��'0E�ȅE�lȒ��P���D��	�����D���7L�̯x�+��r?�OIי�Y>ՙ�Y�W�(�_[��K���%�+a�ʾ�0�A��*���X�~?,o��]wJdI�= ���L����6�y���*�PT$8y�̷��2��7��ͳ�=7[�f�X��	�F�@�+K!�ѣ�(O~��y1ju����F[�I�7�h�{�y�$	�ՙk��d;�d�����g�t���Q4���W���QxS�<�S�P�C�n<c�~y�t`^w۝7~�&�n�s�d{�SG��~Nxg��{��o�k{�sSq�lme��d�N^�4O�_��r��v�Y'������v�5v��+l���q�wmí�V������|���<�j��=6�/.�g;��s��n�Ŷ�g�Vw�����.���MXR���/��=����6}�Uǯ�k��������i�Dck(�������z���e��<qפ���=�>Ǿ��V�6���g��)˩�6�݈��������{��?��%��P� �N `-j��O�1{�ӟ^�S�_�چz���g<���)NP�ϔ��p1�&9����MM�_D~r:p^	HzyV ��O����9�������g���R��\1}�y�W཯}�k���s�W":��������{{I�����l�ƍE���z���dE�J����2Z�N@���￸�'�\���I���A<^�v{�z��x����_����Z��/���j���:�M�2�f�~��V~o�W�s���[��0�y=����@uW���l�p���~�|�@���X_�z{����6�z'K̔f\t�/ߛ୅W�5i��M���Th�ۭ^����� ˻��Ϛ���]����
E[1b6��P�lz|��{ljbk�.̕J�ڻC�v�ZЬ7��w�5'�,��i��qk��b�����6���>n�f'�l5��D��?������s���*\�s�.�I�,^=��������ߪC�^��Wޏ�PU%�}'_���"�*s=\(���x�;�\��)�q��0��ˣ'U}mM����_"� urN(�L�0( ,<S\��_q���(\=^p�siycD���,#��!�2�������jqر{>�$f&�_�I?+!9D�ShAX,��]C*�>�5�8�Ґn8�*�+ml���q���жb;���i�9x:')�,�[�qS�§5��ܹy,���<od��֯��n�޺2Ϝ��M=\�ݙ
����G��T�ߛ7�v�A6Sk���+�v˲=�C;�C;���6³��w2����jZ{��t�U2��� Rs��}�o���V��-�3N��j��
GX�sy�@m0����y��w��X�.����k��h�����b�@�*ǃj)��c]m/��B��&\���{��6vߊ�RXiK���Q4�0��10D -�r6ж�Bǜ�XFn]�/�F���
�,Ϋ� ��oe͗zRY���2")�^�S�D �ǳ�p:�d�^e�@Wg�����+���O���
EUJM
��e��TORCb�����{�\��S���J��4�lfe���m~�:��O�zBsjǬ9�GVpI1�g)��8V ��eΕ&r�ʿ�;�̑ſ#D�UI��i��X���v�q۾+KiX�f��6|i�G��I>f�he �G@7|o�N��j�]u��s�S��vJ�,P��f����\mQ���٘��Z�	Wɉ��-�wN�BCy��B{w�V�@�ffb<[s�[xw��Zs�8�4md�SY5cX��=�+�o�܍H���b$��՗0r}*a�|j=�E�.�9c�����������K���9ʩ�q����N�:7�^����[�R/��Q��P@+V���f�gl�6��p�}���pNK��t�< &�R�)n�|�*�@T>�ܧh,��et'��5q�@<��bw�ب�����,y��(F�Df��}�ӟ�rh���}�|��u<�Z@�vS> %�ac�"@&&�4�&�1���j�Pz�[P��! �\.���gx���V����kc�vۦS6�^��A@͙�i������h�tuѺuV�xӴ�+V[sroXfr���Kt�@3?r]h�c]��ѹTN��z�G�p�͙	�p��lە�<]�~�`�f��N����ϴS:c�X,k�XE�eJU��̪�y����ȷL[���xۺm���7HY�8�y��Y�r�5aw�F۹d���\��N3VY�&����m^�5�mq�B�0( L��k����$�����w�f��'	�s�9�9� ���Yn�@�B2�ɑ^$�`�1�ȍ���j�>�K�7L�B��9LZD�׽�u.�>ң�+�nO�'���N@Yyb���3�=��$�a��M�ƀ��
%�.��M�a\�em�|rEs�G�K,;m �H��H+�Ej�ب����]�EH��6��w�P��~�j�8�@�ik����73=��y%¥��(��c6 ���U8��Uu��&�d:����� �lƹ:�&9L�0M<sp�\����F��wk��;:I�Ɍ��\UaYY��v���ιl�Tr3[hW���iۺ�� ��0�J��S�U�<�i2��'�V|��Ĺ�4p��4z+�_(�"r=�!>p1��  G��z���c���Հ�������� E������J�Wޙ��1ر�����]�h�g�@X[8Ś�*����F!�qx,�����U�ÂE}���������g3_�tG�)���59%�+����p��0���z�D��Ü9�ʐ���.19'Z�a N��)e��@�M������@�,��g>�0.ٟr�W������i�^��X��EV���M}��@��z�_Q��纸T{E���f��1������w�@m�L!���LlN�* �<.��{1���i��Pt��iW��΍���C'��4�S[XT��7��ԖT�Gq:��Q�q�Mz�xZ��s�"ҬV�.�jR�]{w�$���NP��Ұ��Ǆ�~BG��).9�vfe��*�5��\T���`�Gŀ�m��M@	@�ϝ�@���?��u�T�RW*uA( ݣ�7�U�Uq�ɋ_�b����E_.��f�-㍶��H^-NQ����+�K^�9��@[�[�y����P��vh��5[Mw)#H ��8߲+��>�9��2�d۾�R�8A��n�`�,m����)�<��6a~(}�|$�;���(V�(��̵R�^��Rm�9[���&ݭȝ��8[���L{ ���Y��Ľ��sm6�(.@ZX��w�Ez�V�E>_�%�_��fN�u�_��4�r�j��("+�QNtM:ے�Z��mE��e%�2 .@��ʃnM@�`E�F4����'<�	Ex-� P�:C�+���/�#� �D4\�T�1t�	�	�Xd3�����
U �(έ�&1�I��.J�,���R�|��K�����<�*�Lܭ�L[���� Y��.>��5���7����J�	`h{"��e�>���C��3�wH���dt��1IQ�h� <I	�r#m(c�#�u�y"��/��>qP��?�[�r�2��B~���J�>0�:n����L[���L�!�+I��?��S�l������� �@w֟%S9�E��.G�5H�I��e���+#�0(S�÷�N޴iS�y��Ƥl&��j��_.a��e����f|	���c�� �Y�E�8<S@��(D���.��Z ��s�{���s�k�ŹǓM�#����o���z2����Rq�*m��3
Z�D{�Bb�cx�����d ���r����=�5������<��p��@�]w�g�@t��"�U>�2ŋ�L e����G��v�ًE*J���.��|�'�����[:�OZs紥���`���7(%H�|Ģ�q��=�Q� -*�N�D�Ll&8�3��,��B*דs�Cn%���9OE
I����N!�p�Ù\  ��jYi��G8��5��*�^�����.�85�9�G��T����]
����ۓvB_�(�W�1�Ybr�r����G�^��3� Vn���t���s���$��tƒ� �C*$Q�����B<7�qW̄��^y2ĭRf���x/�6���	�X1b�����|�:�[lل�pw���4=_��'���O�MkN�d�	D!�Ggi�>w��r�h�����n�������]�>�P��qėD����$�T"��qHVt�Nʅ���`q0n K�%?��y�qcW�S�e������I'V����0�,�v�����u�O/���B��`L�,Q[оD��� ҹ�m����y�{�[�	@��������=��U�"@G�@��T$���}����Z���~��ŵ�Cq�Dh�lRw�o���N��x������\%C��[o���Rj��,De4;e�0�t/�E���`�߶n�l�ܱ�t��4�$y�>�gZ���=��[��:W�I'�����mG�N�;w���xK�lߠ��Q��Ϯ
b��w�q�sC�)���~O���4��ˤ_��lÝyj$ab^_d�♧��EQp}���΢*R�[tp9J��,$}��~Y���$�W��pT�&���!^B��o}�[��| +>N�#��s�Ҏp�WY���Ec&�+��.+����q�	" � �r��>��'����*0�$#��]@�wڋg�r��E]p�${� 1 -�k�����-��c�&��~������o,lH�Ӣ�C�}���s����s��;��/F�؋Iғ\��>����ݜ����b�x3�=���)��$��=lŽ���f��1�Б�l>3(4VxM��3[޳
�NQ�>L � ��U9d��/���8Y�r,�K%t��c!����c�t�Y	��R}PES)]�Be�>๞u�u��V� 3���

��E�)q]��nG��DP[H���	k1AOyI\�~�wY�c��rn�^`�]�����\pA嶯$.�2 �x�0n	�ϫ�-�I�H��b��p�l������ �R��i��(�M.a*�m1��Q:D�^����(��:׏4I�{T��j�8/�>�5��$������|,�e.%fR��Êt|�(x0�D/���qwYz��,��7Hb7��Ti�-�|f���=8C��z�pH-@�$��ۅXH0*-$j*���&ф�o�~�=���¤��n��P������X(����,�;��D����)3�!W"�B������8j��2�:'�~eC�1�+s��p�1)�#�R�;��+c۹H��#ú�
��k��^j����>pV >����e���R& �Z�?�J�ti�vz��Ń^��
R@���L>���6Y��ۅk��E�:&� 6�.e��y�C:Nރ;ɗJ��]l�6����|�+E�ȟR�v <�e����ܘ�N�W/NV�m�>��gWy�]y�'R^�},$�8��7�3���/���hS��Ё�'��Q�I�����l���Q��Y(�J�Y1i!U��o��T>���/Rw�
yoH��'H�#	B}�����z��p�Ѿ�=L~Y���<KN�;��&͸��@ ������d"�Q����Tb�`E�t�W��e�V�Aؐ���K�����!'�CA�6e���կY�:�8�h�>��伸O%���/�H�G����Y�p"Q(�?}#C�5�\�*u��A��1K�P���&6�b/
����2igE��U��T�%%.����"�8�����z�`��BE#]����<�{여���}:R�ec�ށ�*	y@,��*Ecu�V��Ζ,
�R���g���Iݢ�%�	�۲e�O\|^�?��/��?��+���	�O����7&]`y⡷���X�$&5�� I�c���b&�Ac�&�0P�܈@*��q��2�ɜ�IیǺYq>�*x�� F�������;*��rS*/�\/C��kI6bA�'��\���$�t���������:���o\/à�[){]��8=�2�!�<$E*���K��b����:���or���d��IEh1 �"���$�$�1��ߕ]+FaJ,�m���`9 ;ۗriƱ8jNV�2�h]ό#
�'G.I���-#W̭�D��T���x��X�P,b���E"g-_�����rD�&;��'�rb�Ba��j_7%x����$.p󝅝��uk�@V2�< ��r-����]��w�Ue�m�Hc-�c1��Z�<>1�� [7�	�6)^H�)�Va�qXvLqBE�I�0�>yN]�mz�ݫK�V�yZe׻�L�p�d��؁�%�~�����&ˬ�G��>������c�Zkҗ�{e�;.�gq�R)�f_�M O<�Y+~�L6�xT=d ����BE&M\�b�zo9������'��*��r���M⮝�>3�B�-�V�,�L#��H��
M�&%������7\o�Y�~[�;b9$.VQT$�&2Uֳ���n$D��)��u�_�B7\�n����Qc�~�k����<���7z�BpY?M{t���N]t�����Qgy��y�Ҍ� ���~�"�0"��A$N6^��ʵ_�G,�Jmp(����A�R�,���~�m�ۥa`ҙ�W��,s	I�{|�G�$�
z����4r3I�-$j٠�j���m���] ��[�[��<��f��w"E�.����%���Y��8'8l&x��C�s88@E�<��"}d�h�;u��X̡k�\��s�Er`k62,s2j~�Ї>�If���#Tvc��Da����0�e�}�Ӗ�L����uE��b�]�f����E?��m@[�K�.� @Y|H��+�|�� ����:�z�e���V�*�8��ba�q��v���[�y��5{�]$j�{���e��ܕ�DG�./4��q
Q������2��4o����G�
h+��Ɂ�O+2le����*їg�ʿ������H(&�#��)$�e�b^�E&U��G'�؇3	��ɘ�ݟ�]T~��RVhm.(���ߙ�.���@�뱋�&^� �zI��e餳@��cp�W�q/	�����W�zN��H�� "�b��Cq]h����@�J1�6,v����6�o_��ID\"�1��:�x�V>d� �oC,�&T?R���U�mkn���/Z@(q^;��Gz�� Dh7���>�ޅ������-Y&�."�VEQg�H���pDM��; �,�t,I��J�Dc!bP��	/.�QS\�G�	��u�1X�{ ��p+2�H����9�����ݴ���b�>Y��dH�#�q8X��~�Jy���P��Y�Z�+���Qs�"9����$�d�R*�}�dU�h|�{�͵|�5�&P��8�r��H�f]'��j��_|�}�/ٺ���;��_�UIj���&!����7���A��|j�犸;������P����f�2��~ m�>eEG�A�z����A�Z���� H�M4�+�O+bb�R��⠔`�"^
��)�0��[��0~^��,�Gz�u����98�f�/[��Ɩ<��+&"�~�<��GL;+��|���R}{MB���\*P��e/s��_��>s�z�ܭ�����X[v��_R��%j��o��|�<����X��x��b�o���d���-!&a���"$���6�v�K5|���63�SŊ�j�C�����un�Vq�,YH�Hۿq��"�\��� 
@h��R����߉�!w*�;q*�a��Xp����8'j�j�W��b��JM�bB=�<���{��mo�m�1��v:��p��tG������9���˂�h���	#?�2�^V���jEj�اt�	thg��[�y�L=�^���7��ᡂIPgP�E1�_���`����k��4F�e6C�b<�x/,5�[\�)��x�:��8��.*v~q�l�I%RԲD6����O+[�6I��	�%]�����9�*��(�&�RÁ���8��nK0���̳�Ǒ]���J��@��X3�� ������dIF&�b1j�7�me��9>�;�p�yp�������=��ݨb�3��-��dG ��r1������%dV\^��+���x�+
���LZ�;\�s��]ФWe��^!�'�(�eY*��W����� �8堒�#&�n����084T+��� 	��4q9p1aR��J��� "� ��:3\q b���@��G��#,�<K�)ę���Q'`|�, ��z@���L>�M�I�� 8�K(7 E���5�V�5Y�eG{��%@]h���W@�>%Yl�r��(5m ����W�@�k��>ش?�xy@
�┕�O�y�R����T)�﷜���!�祤�C~��G���֥WU�(��R��{���A@�\Z\ �?�k0���W����ɡ��E@����XZeU�	����[�E�8�^`���;�R�Q�<���W^�X��5��r�҄�w��R�}|��?9��	��!��X܎AZ�U��3nGk�#���@E}(*�]�]ғn�
8��mY�<�o.ƙ�O��.�d��l��&ڲڊ}�K��o߾Ӎ9p�d��@�C~��2,�|'W�\�����rP�g��*�\�0�ɑЅ�dE��D�� e1�l\�Vk7�m@�G��ll�s,�e6 ��
�p۷c��̳Ͼ_��7u����\�bc�����-���3~W�YR.���eQO�Y"s�@R��XT�T�H#�m���f��+h$��/��ڽ�@�k<^��H�K���jҲ��O&�NR7���2pE�crx��<�x�ø������W���0�-����Y܎&�ܨ��J�z9�kwTY^нD�	�⾬���/��Ѭ,�Y@"C�ʬ�R�W�uYu׮� �O~�E����Jܢ����x�
��D-���7-X���S�ԩ��Z��w9�����X�N�>C�sTHŲP&��Eⲩ�t�
s��Vm�l�3lAKQ���Zʳ���7ٯ��f�K=���]֚��n��#���R���h���Fi��v�?r�9Yҫ��]⩩,+~��E��Ty��#���k��;�HH����B��� �f>C��K4drQ^� -j��UF�	Ƞ$W)|���3��L��+P�:Ĝ��:�-VsvF ��bƝ^ܔ8Yލ7�wY��F;��F�K�|@e�����pc��S*�X�G:���p��-ݫ��Ny㭾e���W�¹n�Ρ�� �s�6l�͎�� y��O����=I'��F�Y�W9�}@�#|�sf��%�D$Y�����/bX���|��xK�^ɧQCp/\kLd�R(#��xR�9��^��Ke R΄X��w)PReMR�ʊߗ�O���x���/u#�$���1���$,�q�3�<g�ܹ�&|�z��dW�_Yĥ���x;��^`�@0�rHb6m�w��K8P���+�B˽6M�g����O-p��/���I(�"_n�#h��������-�]a�f��:�DO����N%g&��m �t�_lLG1�2!�C(����ۿ)"�`�п
l���f Y�@���LpM��ƍ]-����=�b���+������g�{Y}2t�Å��E���s�e��\�3>�Y�$�����Wx�}��j�'g�;A���p����l\�2�	x�w^Y� ����&�ZL���
����X���?�A_4�԰.7��~����N�P�b?�L�\�n�C.Z�-N�G�A��Ŗ�uΝ��c����l86�Z$�Q�ÔPVj
�q���P�p��y���u����]����Z�h����U[�Ĝ(���� W:��p+��h(���� ���:�`�����J��H��qx�8q��9Z�����]I7vY���{�TV8�k�[Β߫~s�����Hb��3\�Ԣ���X# ^
0�F��2c����)_}��]7��Q�I��P_*a��vwWQ1V݃)
UI7�u:$NZ��LT�XN榰�p��=�Z��ٰ`V�^�����܍#Kg��Y�|��쪟_�V��uY�i���q���`��!	G�� ܲ����1�X�����p#�|.N����|/�)��2��$#�R,��s,�����],-�=qi}���� )o��=�t���Ǳ~!Z��'���?����݀��t�e�3�
=0��XD���P�rd������gjCD-��,p�ݲ$�U��~��Mvh�:�K%��D�M�<R� �}�ؼ�[�M�4`͸��K�m+ˤ�Kǰt�}ʔկ�dyA.�߉�t��AY�D�9��]�.ʍv�ҥ.^�Z�����4���/��2a��{��<cW�����
[�ˤ�,L �fܺ�`�D�˂���)�����Q|����(%%���&�9GhY�������V�?ʻ�Be����	<ʉt��/�.��EkA����%��S��?�_����G^-���?`�r� _�����"z�vr�0���Xm�<���$_��z4[3��n��4tɶ	ϗ��J!�5G�Ī���_���<�@` O;K�ӏ�c�qΥ�.͞�0���%�o'���s*�J�vS���P���&���i�<6��4_��r�̧$[G�Z��' n�kO�㵒Z�%��a<uL[]�����H�H��Xj�gJ�J�U2��e/�~ǎ��9�Q��Q(V��J���k����v�0�y[ҰmnC`�ݖuZ�t�����=\�~7����96�KSL��'�WQ�9i�������8a%�V,��� P��������vᯌe���8�j�f3�5M��(��%���Q���9:?I�j����rs�U��Yd�d�`��U���l*�y���� A�������@��������8�+�Ց>q���7���g|j�f&3��?w��|F��ejc�{^��4Y�:�x]��t��礓��O:��^�������?����G1d�b�������k���o9��~z�/����LX ��ڮ��^e�n[��8�)�V	c:Վ"I�63�(���hA\	�Z�ts��Yl*Fjj�l�;���� a �p �I���;F�|	�Vc�f��ÛB9��5�"�nR�𢙖?ϙ�*�7K���4eZ�u;�V�P�Զ�����lێ�7U$L/�r0G��T��<�87�8@	��Eo�� O�^nM�*��V�Zr������Ėr��g*��!:@�	�;�c�؍U�u��_��b)���}��-���=��%y_9���[���ҳcgy(S�@��0�j�����h#g�:���w�t���pr���ؙ�V"�?�C��&�)����BZ�e>��d��-����� ��-gR`�����t���:��[�����X3 W�W��j�-۳s��������U�Z^��J���~|�J�:�p�E��=6���g�P��&�w���G�K[�]�Q#PlkU����� ��Z�n�O̴�|�РM�:6���I�����}l�e������HN�-��4���q��;�#�dѫz2=�h �bP�U�s�Y�Y��$W"f>�L<�,z�A ���w ��F�#Q�6��Kٌ1&���#��BIV䗬����ʿ����*)���c�.Em���a�J�C�-����(6zԾq���v�(g����X���TXv8X��+�����q�]vL���=� @a�;P�$�$���伀i5�y�9Y�l�(�N�v�c�u~_�fS�����lO �����x���ٵ�^�}�wl���#�����9�16~���]�'�-i:��`>ᔭ\��������jm #^�F;�<L;̟403�/��Wa�]Ͽg���g�'�3���WM���Ya��k���,�f�>�� )$�����F��]r�#)/�ַ�Ҽwbܹ �5��U~��f1�m̭��K�c��\�Cg�j\�/����i������W]u�'�&��6��]��ꖤk�>t���s�t���۝������\��Iunx�@�;�8T_%�'�=ȴ����B�W��8�-��ra��zRw�
��M�����?Ӫ#��G���Z[�g����\�+���A����[?u\�F��憦���9w�i֬ݨ��Wn�z�f*#v��g��g=����Z����'>f���e���o�/|��v�~��{�F�Ks�:7��::6T�m�۾f����W���0�ø9b+���s_���>p���	�g�6�����A��<�iV�v���m�i'lz�M����m<�֬?��Ҵ��SN:�Z�G���S�<�j'?4�a(+��g7�k �?��������+����l�5���q�6���OcB�=�rY�I�5��
�eƪ&&����zի<�8����Ӊ�5��
������,�z�K��<\p��S�gڲ$�DQ�b z�ސe�T��=T�ʢŁ�"fLx��%�^i����Mѓ�.Խ15m�{���E�l��;�f-�<)��N�����'6����m��&;����v���~�FOaz�}�@p�>׷w���`
�9��N�Y�Fs��|�~�6kOWl�nt��c\�*p����cΰ�Κ�8UbvmC8.���I6���m��Xܲ��?��v����v[������w�Cl�����yn�S�z�����\�%K��v�S�����/7�E'H�g?�&n��:���S���i�[�-6�s�����T�\�3Y�g�?�yf{��d�2;y�j���P�����Y9�ɜ��s��/�3ϸ�;�cѯ׻"|�Ɏ�3>�$�AO��y@d!G<�%� t��%�(���Z�g���X�Aʒ.q^�:��w�;M�}�s=����L���ώ_��WK 7���+�K��屯�d�Z����>�IOr�!��t�JCI[�O�u,�,�Q.�Y ��B�}FH7�*�-&���	�1�);ǦM�
��xj|bN��^��H��o��A$NG��|La|jW�mǞQ���c��=����dbyn��ڭ�݃������J�>�NM���Tmzj&�MŶl�
?���� ��a����=Φ�U�L�X�Q<-
Ǌ�tE+�tʕ؅j�����9yȎ�O`��Z�ʶ���c����c帇ۆ�և����9��ǙM���㎷�c�vփN	�k��N����zV��?�����}Rxo�w�;i�j;f�	�Y�s.��뤹*����L聳�<˽�����w����.�r��ye���g9 Kle�d�Fb�	���x L�C�4�7�8V&p��C
�&�2�r�&*�={vۍ7�P�!s�n[�h�m��rq�~���͍�U����*W������	HӾ,VR[,D�ő�Z���@�q�������7��K�po�4�{��e�NHp�e78~gQ��8��6�H��1ȶf��Y�+�QAi ��m��������Vj����>���h����;,x}%� ��v�����)�s~�n�x�������ve�l����,T�m���m��+�`�l%眱��=���^��m�x���V>�֯��qF���v���	��]����O��f����|f�%Q���'���΍�;�>��x8�N�v����N��'E;��P�.
zL�H�Y�ֹ�b Y���B,H_��9���P~���ܸ��C��7�1���'U`,:���ߑ�#���W6��>��Yv�)gugɗ2��*Y	� �� a�
�*97�b��W
f^ٵJ�@��w(��؏v_�,y
���E؅r��ՌD>i�iU��aUl6&s.�n#�C^�أ")\u�,���(��x�BDR�J�]�?��,ڮ.��v7��j�[0��V�L�z,&������r�Y���j�{�Z��&Z��p���u�����?P�Z�o�����ӟ�f��c�h���n��X`���X��C������C�H��ߎ
��y]\e��.M��5gx�r׳zvqR��������g4<����̴�:P���Q���g�
?�^FΚ�����1�1����s�ٺc����L����Wˬ�:��>Up�p�p#���қ'Tр w, �p?�Qe�W
:E_�׀g|�ӟ�rq�ܥ���\�b�wQ�"q�a��}a�Jm���g�lgf��^���70��O�D�N\v��P�Q�Y��G=�1v���n���qXrx��0�=�!��?����y�s��ٛ�c�1�a|�>�)��ھw��M#&�@"Gj�wς�E� �����'$�Im'�ю�2�x ��2̗����) >�*J�|��0G��e�d�A�N��N���$��m�w�t2j��5���t�#C�i��w���dq�ֿ��'��kw���:�j=�m��I�d;������ss+I&Z,Ҽ��2?���Jc�TI���ߚ�'����fA� v�d��W�y�s�[KP��Ts�Re���� 0�3P�*�U��m2��
 ��]҃�⋡��$Q[9��o7n,Bu���L:�h�nr�Wn<��N9��'MaoI�7���챏yd69=\8��~�����n���s�8�j��9��{YhY���zev�7�a���rGٹz�s:x�h��_Y7�1,^�C�◾�'[���$�}��m_�v���H>��m�tw��s��=�������~að܋D�<����7� ���I�z�@\��x{ǻ>`ër��y��c���/�K��=b+gFZ8S���rN����ٲq��im9I��H��g�ou�OI�$GT���3M�;a�7o���p�u�R8O<F.%�#=@�!�E��e�eP`����,� '`�
����s28�c��73� ��{�61�-v�`'�&311R�v��f�v�e۶�f3A�ƕ���f�|��.uEu��;O���C��PjT5p�D��޽���Tb���n����rk��[�]���lf]��ZG�7Y-��Ֆ8��/W�Z5ۏ�����h ޲_8�(E�@&���#�D\���@q�%>��u���A��M�I-�U^�Bߊ�Y�����׵,�0G��0�s$����vA%3��G9�~pqT�� ��yVHq�j�h�9����z|fB�� ��[�X����Xh�E�%�xY�j �J��\�(�,���c�K}��v�a�U�q$,"��&���V������T�'��7u8�J&���Sג�qNv*,2}���{#�h�`M ٝ�p�q�E-���~r��P_�B�����8��]�5[���+Q��&��ơR����\��tD��p�%}���|����R7\؎x�,&����;�V�n��>򑏸�
�I��W�V�Aj2ЩJlJt���]i━��c��<[�-T n��ب�����}a�V�}R�w<B$q�x+��:3�b�$\�O�a��d�*�S��}�z� �7(�ܴcj|M�����L�4ds�]��rm%J�q8�W���J��������)��D�kN�R����tX$����ɶ6�5 +��Cj;�ڃ���݉-d!�E.L�</�p��/�؏+���E����Y�*q�����^�� =p-��t>���( �>��w����^�7#0��`Ubm�(��tc�����@c:Zy�~���D�-m���t�t�����T���8�f�Ԭ9G�9e7r�kղm�;��Z~mr��*�"E�e�}������\���/nZJ����N�����.���h"�������'O?bi� K�����#r�X&y0�'>�)w"��kх�D,%�3) 7@M�� ��B@�,��$3*����K��a���`y"h�-�w9��W����BKa��"�P����4OzQI3pr.��{���V�V<<�)�L���ݯI��\���a����)KMw�n硍˜
*�w��>>�m�A��~��s�C���/���8�/��?�)O9�:�厂���G�5�A���*�e���b+�G�嵑��d��w�,�Bڵ��N����/~������GF��s�#���xD�+�C ��hA� ~��Dl�c��x���@@$��8W�e�y2�0`P] �RUh��o�����*�͝�(���+U������3���Oɜ���]K�w����{-e��	�g�'�Ci��K"�DڝG��=fE�Șp�@X_;JH���d{p1>p�S�W���\���9|�|�1�d`:���i�n�ߵe��"e���PH~�e��9e�Ad�0��?�G	'�d����;�>���9�f�͎���Ϯ��.��w\�C$�_62�s�|W/��"��V�Z� :���z�x!%?<9��2�n��c�s�Ez��q��n��F��(#�>�j��u�����b��	~|��E���Ks�f%�qΦ}��<bbO$O��z��,93��8a'i��S�wǋ9��O�5�|Ձ@Q�P����P�m�w���E4��4�ab��z8_$0�2�z�ʴ���*����3�/f���e�C��|���#��\Q�_��;ش�,aU���E}�����~c.�K�\�; ��瘞o>&~���N:�D�ѳ��/-�pKK|�s��!⩕4p���C��)�	c�����w����;��8�*���^�qb;q�F!$M�TT�(�D�Th$��!�sH$��SP#E	�"E�8p!U� R)"U/HPqDЦGD���P�FM�رw����w������ƻ�y��ݝ��ٙ�}���}��;^�N�<r��4����Q���S~VǶ����[Di�����?O_�-.�{:���K��6>Ts�=�Vj�P�#؈Ga@�LS�n%����j�O�%ܫ�dU�r;��J�oM�`�On�+�cb����8k���s��[P�X�dUl�Kk�d�c]{��`���c*y�TT*V�H-f����H�n�������*�'�?^��^�'�`��ؓagg�����GI�� !z���z�~�;�ڂ�� BV��R�Њ�zj�
�%5=�^L�h�,sb��N.�m�&TV��.^VΚ>�Ulio�h&&g�W�ɽ��+	�.��:���_7��7�4�ݾNk������>y�(���4��߽�}��G����y^��~�v�jiG�((xy�@^{�(6�u�ie� #�.�pW���&2�㑷�ET��c��)d� ��d{��6�y�~� AiX���=p�43n4	l�Z�������@�K�� �c�A��nZ��>x���W@�שƉ�(N
y��ѯ%�cQMu�$���u��k<V�M�)����l� ���뛜v_��s�/��f���-w�wM����A�R�z��ܨ�$�}�)��g�s3�$Im8��U&&��t\SFvS��4���bhL�,`]�|��{�~�Gͽ�G;7�����lP��i�Z�)m� ѕ+W��cߍ8v��	��LY��9���J�s�mc��YX�*SU��]V��j�Q��z���lU'La�y��_�e@�Y�(����6�"� �8���!�P��kb��|���_�U��o|���׿M@�O^|�y^�{��ϧ2�W�ޓ��X�wئ�-���T䅀P[��������O�VW��R=� �����~9��ۯ˧Ezoa�PE#����g߹c>�T��]�fr�T	�<�@v��Y{��t�;v���ՑB)-�ܻ�w���U�$�s�&A&�ĥ�?n8��/�	XE\�۷o�m�6�,�t��|n���ԋ�\	�(aU;U�`��5̅��@'&��$���5Z.[Yf�08u����Z�qZL���������h�� ��r��m:H��Pdc&�2��~��{�ͫ�~2�m�:iE|���i�jy�.�0��j@Q�)�k�wz�̙������-�|�����-' ����L�J5p�Ec�����hI�����������*7���b��̞��ћW���m��2G��W���]�$n\� �N�[�Z�f�D�
g,�\$.Bc�clM���A�M��g@ij� G �V��Ծ��Z��D�=A�M!�:���u��N���̬��t[g�%�l�ū�;9�]�M�LV) ��Z|ViX��j�UE
�L�0�x��}PZK1�8�k��Y�S��e6F���	_�x�"�$ �СCɽ�SGx����$yQ��}��>a3�%���6��a���^��E����z4�X��D�`5������d�}���L5�a���fֆ<^��Ax9��O�8��m�B��~?X�jh+�ܐ�>�d����l���VX�V�B��I�F׀׸��Lx����g�Sa)'���rYՃo���}�ZК���QZ�J]��ˮ����z�D3�#�0��Ġhˍ�?x��M&W�D�-���|�ޚ�y�͐�?�eV�WC�v|����;ʓ�������Lx�.<���j����#���s���.$߳l��ɓ'������X��Z�|�gݻ��%�|��h�oQ��7G�����NJ�C��u��e������4+�	�|��o���{i$ ��F�巿���؊�A�]��""ҭ��*�*�o���H�5�M�_>Ud����fM�\M�ax�}h������*k�!�_�u|���<�DVϿ��[B۹6��|n��߽+y���{:�l��`�z?��!-)�¤G��Y�S̨M꧍h�R2��0 t)����A�R��	�\���[��=��A��U��`����Y O�,��ҩ� "�TX�G��*]�� �n�2:\��2<�7n��^��5l�u*9&R.���%:��X�-�:%���%��;���Y5�^T��#vf����<U0�ɖEIi��*/>�G9\,�k�d[Y�����B��@^�p�6-�%Ao�0e�Kd�hS���E���_���>?�=�N����?n�2���6�nI�&�E��ԛ�yRnY�<x\�uҖ|��Y��;o����L�G�����{u���G��)��gp����r5�Q�mKҜ6�`��|�(�٢d�F:J���;_���5�����������Z��G��v �me�~�ײ��&��ۥA+�"��������������x���j7��������A��>�;��τ�&,�3*��57�i���ո`1�O�3jV�h�����V�uaM2�{�*\�,��]@h+�V�l˃d�(�k+��`��Kv�-�M�+�s#V����{	�L��<�Nt)m��e�C@��A�fg�Z+g�c�R�#���u&�]�w��4��(�5�)M�Z���&�D*QL�Ut!�?$�{k��C�s�������W�H�&,���L� O^b/J���b�T��v����_)׾���61>�:u�=�A�$K$;1Ysq��M��I��[�(Y� �Ǫ�ro*P(Y�`��:�q {b���n��[s<��&,��3,�y�p�;1	�p^�P��4��@C,�*�:ڦ��PB�m� &@e�E'E�Z�f�eї5�h�uǻ��@��+��
H���I`�ASzeL��nC�Vǧ��ڜ=�ߓk;�;�v싲�����~<�2��Q�߳�$�"����C
iꔁ�:��E���Ͷf�]E�꣩;	��͛7�{��s�`��"E\K�[ĥP�g�#Ӊ�4] o��f4 U�ˢH1Ük^D�l�,}�ۿ�S��=o ���O�m����u�Q�,��R�7N�!�Ə�a�o�~c��9�g�H�0<�����nsm&�f����l6jY5a��u����d�S�s��w��iw���lܫ_�K?6�徊Lx�3|�WYg��� ��#�BF���xP��X�ɖ��4!�{0��$Bi���[RC�ݱ�S�o�e��~W҆d�8�u�ܩX-F�LEٙt�7�h�W��Q�n����]Tz�{���
bp��"��{(T��ls��e-���A�I�Ԩ�I� [ړ�҆ݓ����� ��9�{�ާ�[�F���tQB���Q�����:�m�Yj�� �)��N8Û�Q��,� T*iO ��S�y�|&?��J@_�g��Q0YQ�Ba�QJ<W�[�{�X�U���T��.P:�^���TM�c�"]Y�Ԭ �!}+o$��se�m6�D�.hf�j����ݤ�����`M�)*Ǿ��ј�e����;w�f!���`4�
d���
d[Z����1�e�a��yev�@v�-�@���:Gȶ�^��k��o�[��xe+    IEND�B`�PK   |G�XEm��O �� /   images/f99a6fc2-4a50-4dfe-be0a-52d397e863dc.jpg�w\ݺ6<H� ��4)ҤH�$H/�Gi�A@C�&����t"�"5
қ��P�����s�{�{�~߽�����Cf��*�}��5�֐����sPUuU�� ���4<hNRQS��������9u����3g9���Yy�xy/q]��/,#�YR��E1qIYyEEE>�[�7Te�+ʓQQQ�R�2��2
������G������x��d��d�6�,���d�}�?>d'�)(���О:� #'?AANIIA�	����$n�dԵ��qe�|����Vy3���&���ZV��������e����+ܾQU���704���Z�<���wpt�������}��9*>!1�erʫԬ�ܼ��¢���U�kj�ZZ��;:��{��GF�_������/,.�X^�mm�����������_�C��9կ�����������I���TV��<�O��nŽ-o����d~�6@��'=Ï�դ�Z��kP��Q��֠���4�&'��P6W��Ǧ�"<U�$�="$����|�VS�bE%�6i��QH���Ϗ�v��)���v������W��	�ŪZ(�d&es�����g��@�.��P|`��v�z4T��������t�YU"�~�;P��y%ݒ3lE����9��;Q��oS��1���..^V&X�-��I��3 ?��J&�`��d��c��is�w��D�5����2B�P^C�C��A�Ш<d��g҅ L�J�P���B	Y�$�c�ׯ�:���N�B��r��t� L��o�������`�K�{����
ye�V����zӇ�7�Y��B7.��>��{�淲�;'U1�m�x��G��4:��;�������@X��#�P孄�Q=>�@�Jň�Q�o8r߱��*}ut~�v�8�H���z���(%��êw����&����OC|��-����R�ָ{6;�26��H��K~�S���J&:��#�(��+Od��|'���7du����Gh�j	�i �ڐ���ɡ�A&�[�����dlM��&+x�֢����*����s�J��ӫjLT8��ߟ?�t��p���iYZ���G��*�uǂ��0�e�^a�4���P�G�_��u�T+.}�3��󁡊�c�Uc�'��{���Dŕ��.}7�@U ��c�w|h�l�����O&�}h)�^H��>��4M���J�	�w�c�a��Pهq�����[����&��e3\{��4y�s]�\I0��J��h!������wi�dnV�q	���z���p�����{�Rd����q��D�<�<����'ǘ��<�X���m�e�8�01�ɯ��U��]���6�����ӣ8ǫړ̞4!��1����֙��Ǥ���sW^�w�t�*y�L��	��!��}p"{�v�\�`���ꪸ�H���#"��u�W���"Ӄ����Yc�^�g��j-��R}-0��M0h���(]�iV"�SqCg3���@���~�*�s�k�M�*`p��`��3�;�pM�k�s����L!b$?�>�{wF��
'].��ˇ}S���y���a$�pf��ʑ����!����{�B�"�⻈���o�,w�x��-Z�����R�b����:e��Nі��S6�]ܓ���nks
W	J'�3���.b�6�$P�
�`٭���7OV����v��s���݊��;{�Y������jYw�9`�l��HHg����[T���*�í��-c�+|3˾Yq�e�T�^�n�V��y8	����uu���%Q��-�BH�&�����v����Suk_�ʢ۪�U~T�xB���n;���=P�k�a%4�>
]�2�3�� O�O�&���a�ht��4|L�����!��x���lT��+��쇾�a��'t�\�`���4�c+k�r��}�>*K9\�3*�cN㑱.����K�܇���͘ĺQ�~_%td����oL�������us�7����{�ѓs�O�d^�S{�(9y���8�kW��)<b�gj�㭧S�+���mSGY�U��p)�չp۰���-ט�c���9h���fS�萯yw����'�	�2�MB6ɾ��g0�9�QџKO�ħ��� ��}l��R!����I��)�l��A&΁[։V���ݻ+Ji�3��w&?�	~Bm;��]7����aJ��&����!���{�^�`��XM���ջC��-Mw�	�9�HEЫu�p7�5unyթA84�����K;�Q��P�B�B�ƹ���W?|Dn��?�J��M���1��>��Yb���e���hd���٭ؑ>��sN,$���ÀI���X�璔.�U���/�ҏr�^��|�[�7�g�+����^�%)K����e;�i�z���i�ljtx�}1_y�S~�����~x��|�9�d�}#Bv�p��g�gRMr��nuR�ڼ����C^%��>�Ө�:,��.&�Tx�'���\n@�K��l�}ߖ�k��Ժ�J��é^ ������Lΐwl�3��g,�v�śV�I��η�_6asq{�2A	)�3�I��k>A���KJ��s�uo,��7X�E�7�A�4�D�Suȓm�%��/f�3F����g�D��S��'"�����Tj#pS+i[��Zd�J[���EF1��X���o}#�Cq�����D�٠I\���>T˯~f�HńK;T�=8%1�X�p�K���G�L�a�F��[3*H2`�'z-��'k���tိ�����U��c��O�,�M��V'���]���zXL��(�Q�Vv}C�����^�1�v��9tG�]�m��{����A���E+�{�}pԅ�TÄ+��	[�s������e�@���x��l@mJ�i��R�x~�N��s�RO,ނٟ��w6p�<��o�v	m��y��?}���h*rw��^ ��]ݓ����W�
���G��09G��1��42�@	��Ɵ��(�a֐�S��QOj�K�\�\-���"��lS����l'w9�l�=�ǻߪ�~��X2u����Ī�2���Z�s#����k2��QWm��.�]#U� ��	�G��	���u�/N93G�;G�i(ڏ�9y��_øc�_ͷ+���G�ZJ��6��z"k,b�@�̔^\��|[:�^W�ᛙ�?�1ky`��f��.�N�,ϝ�д�U��~7�zxb���M�qȣ�m�T��h��^w�����8m��7(,�nw�1.���(B��{��L���U0�#(ǟ�ּ������7B�%�[�� �]�Dc��<ne�UfN�u�|�W	S�0X%N����}��|��W�S.�ڪU2}L#�t5�+�ZL��O6��L��.d��t�ye������RZ�!���ގd��k�\OQή�R��{���C��t�2u]���Μ��f�T')h���Lw��po]1'X���gS[
����M��z&{�	M���� i#L�p���h�?�to��	�&�=Yt�%�d܂��[��Am7�[!WEڳ�@�+b����l�.H���Q��\Xjw��g�'�ľ�Y����g�Ô�K�����Tԥ}�xv6{�EY_o\��g�|a��ұqQ��&{�N~�������.'�D"�]�ʣx�f���dѡ�ɨ��(J��j�h�|m5<�Ү�bV��Vɾ
���$����H�*I��V?��U�Vc�mC$ 8�#�i��,C�C\��i!�/g}�R�*���l���~� 7�����[
�s	�W���QW��#O��,�Wl�P�OM�\��0����;:W���5�]�R����"�c3�!���s�wE����2�QO5"�Y�S�
)�r6���'ag�]Ɛ�������_�E�����h^�U%ӏh5�+p�~�qb��yr�4����Ne<e��×��.:�e�n������~z�Q���:��U�&+]'������}��`ΑQ�0q�@�r��V��⫎��'�m�oXP���"��o��NKY�#��[)��ߟ�өP�ޓF�8{��ŽAې��6�]lަ�v?T��#�8�t���/�P>T������u>P�i}�a�݉�2��5ժ�KWL�4�}�PZ��-N����ȭo��)ܧ����t�Wj���=/O���>R�I��۱�?_�w�-WU�ɡvlO�<1W�!6?i��Up�pP|���$wG�ǑvE�c���H�b�
�J�[�=��u5�݂���c��AZ��2[���Qm�9Wm�"z����#{�ua�9l����o�F�F�8��¯�fga�ng���3 �`�DU�W6ޙ�X�a,I3�)��-=���{�L�m#�HX۲��g�a��/O
	f5Mp��"��ˆ�#�j��9����<�?g� _�.�0�Y�a�.�G}�Mto'ss�p<�����*�"p}4�aG	pF�TF�(J?*U;��G�/q,(���p���B�um4����T�D��ZR�*}�2Vm��ik�OY#ҁ��F��>ƙڣ;�w��y^����J$��/�(�2'��>����
m�&�U*��u$�}��DXU�+��x��{��pъӧ�q_;:!����9~K��ɦ��"-�G���h�I�H�	��M�P��Ŧ�����`G��qw`��ɻ4\/b3N<�!�(%g7܌U4�ğ^����[�i��z�u��΢1(�/j�q���/Uvۆ���U&�`b�4an���W67����nFN<N���+��FZ|g�L�n���)>��$�tZh��!��)�7�Y/_�ǚ��`գ��{�\ ��!n̻i�!>�ui\�m�U�T������H����v�U�^e�V�i�[X�J�I��kףs�]�B�?R����z�����볛s|���T)S��A �pDe�t��ٴqt�����'��F�i��t����b�H�&	(/���y}�uR�V�%�H�j*�&u�(��ZU9�4�Dμ1Ͻ%����6g=�6���M=jt^���jc����6z�dK�:3�M�����v^�Y�zPv}n�7������u�b}�BiL��1�KCow�5.�~T��k��s#m��� @�����V�w;h3jH8m�>~m�7�( �A'0q�k/��E�D��D
�0�(u��K�տR��v+k,U��#�8� �Ώ��K��G�H �WN�6�.�����Y��M3W<"�,
GəJ$���l�z`�o{\H@\ˏVT��߲����A:
�~f��ȏqfܛe��A�V����-{C�Y�2!��xe�~&w�%����%Ÿ��a�l�ڦ\��
}�޷��X��JR3j�%�2k��/ e�s1�g����6�������o��Gz,կ><4���=�=˟41��RU^'����ݨ�Nkg:���,]zE0�m�{�3OeM,�}�ѝ��� +��d��P�Q[��^Q��K�旔}w��ATFv]��9y�ܡ~J�Kϭ1ڻF��h5\RZ� ��Np-K���!K.wT�"1�v��ck��`�Y��v#@{hFd�D �Fk�Q�����{�'qZò�*�ŧ�&k(�+�b��(� ��sJ0�bY��d����H�Fȭ���v���b��*x���-�u���p�a�Q̨e�h�oN�� �C�\�|��qL��,�$�#F��װ0�C7dه�YMg������ڠ[�`��q�xL���uP�fcFha25cֿ}�t�'uw;��|��C��"D��z�h���;>��&��2si^����e��_��,έ�xw4l#'�?��nѹ�#�dx����Q����[�	�`���||�&�9���ٻF�$���y��S�@P(n���lAҬ�m�x^r��Iq���*bfb^~�e��+{�2]uxG�i����ᅹ���h���`Srh�X�ۧ��Cu���$��^E����ǋ��Wr�P�GUf���� -#oM�k��)��|�l���څ�����Ж�ٯ_J�ӱ-�;p�6�?M�S�| {G��,��t�̯��=Pq�E��$|٫2�Q���<�2o\z��7=f�cDe�ԯ�c��r��W����SF�p.��y@�Co>p7Ѕ����2R��LY�߾jx��3L�2����(S�k�]H,��6��Ď�AQ��F����(�����oC+1m<�σS^~2P�¨g(,x��
�(�YHp� ^F�[0Y�(u ��)Q�y���`x�a�ϵS��{��IT*T�$85k��K|,)QH�����
U�aMe0'��m	E���1�Kdؗ4嫂�;��#��.���r�T�l _(��>�/�Sv+Q^���S��̊-�B�9L��W����|S�����G����Я����?�M�Xfm����Ow�f�r�����r�P��������+-T��W�9�h7f�up̾��Yc��gl� �?���^`��]�.����d����T_�Yu�HbM�p�)��+'ag��cI ��� jS�_��RG#��f����/�����T������1�y��9W:�g�v{�mq���u!nL�=���<K/�Np��M����%�\�Ͱy��pdʆ�����<�b-�;����$`J�������qgY�	 �-gn�6���\�9Q�,�
QF�$���%�Y��R����0��p9x%����U7�{M�������C�[�r�*��.��O�l��\�h��y�15#�>����N�v���.>��V����3a��\�"��]jʫ�|BQ�\��d���JCz%�`z^���b�Du����� 	���'bm��>��g�Ag���$�9�r�8"�LH�
�!Sn�+�}F��"� �g�7�"�L�����E2�y�Ww�q-���4̮24f�!A�ņ�9�S��z����&�(�yC�� �q:\�F'��� �����9�'����ȩ���������O�-r��S�	 �gZ���f�2��ת�����q��EHXZ�����W��5yF�%��#K����xd�a�+�l��w��;fz�����V���9���֤�EL�i�	<�ζq�����$�-�#��71{�QApҎe��#`���D�%{36,��]�v��|3�%BX5ۥu�W=	@)D�`�,�g�|+#��zMه`.Yr��ӂM�3=�{�񱅿q��ן��Y��?�X�X�VĘ=K
�2�](/�K��Z�p(Ϻ����4�!��ɴz���ao�/�5�C�p��i�Ȑ�����ܻ%��'��=q%jm�S ��p�,v����aC��wL	��[ǧR��EL
�z��!���Ϳk|9fx��#ʶ�u�F9;�;�WjO��}:H�#�q������5��jq�����g��PvhY��3!�����Vx5�d�<�?�3XGI�iojf[�]�>	�x��p$��?��R�mn��� Ф��rZi�e��`�ǦL��'�lvB�U���ݥ�rG���Sϧ�n�������o���}�E��x�G��7���n���և�ho���1��1d�k�g��7|uk���tIk�2�%�����=�V��5�}��.���O�ҠJ##���Zu���j���7y9�,����;V����caxrÝ������+���`^	0S�3.���B�i��f%�Vq��$�;?�r��@hI�j�1l�9��qv�ˊ��]�W����ay�Rӳ+�r�:@h� �A[�:�Z�'xk��F��z�� $8�Q�K��Jm�E���*T��}G2�e��^qkM2$�v�XS�Qz\t:�h�x��E�!�F6 ;byq �d��s/�� A����#a*\�;ˉ������ǎ��/\K�*�n⾅E�`}��D���jZ9��6=M5~TԾ��d������q	o�'FD}����꠶��-d3�!L�і���B��ᙗ�/�M�AoI`=�p��`Cv�X�UZ��/�@v�9���lpڭL�G7�Q,2��&߻)�z�\��������g�f�2�v�E	�|��/
(`Z:K/�\���g��@��`�XK ��0n� �U�*�	�c��I2�����P��,�����O|�iv���:߳sQ���`����P�R��?M����G�t��gM�dyiFS|����(���yqn�M_�������0�L�_�U�ϱ:�^O�O���ɒ�CD洂��:�L��_�Q��˓O�*��a�MC!��13��|9}�㛿e�*0;�*'�6(_;5��2�����%_6�ɖb����o1=� �a��s�₥��:ԏ�_\� ;��	���?���KeU{�����Miu�w�.&��L ��7op9�|��I���C*���D:d׶q�%��t��X�����.�]��4��~��xL���y*\�:ɳ�z�95�˯��~"]��Z��-펅�:>9��ГǻK�=�ijG.�p�d��!�E|~��W���P&�wUfJ$�z��@��)�����
w��Ӄā{�Z�l5��0�;����%���=;oF�U5m�I4=>7�j�����K`�*�-wM��(j�K�S�R��A���UYS;L8;[���MM��a�Ȕ����c��pib`��a��!��Q�p���5�_5U+S�
�:qr���26A���!L����!�!���s&��K����v�;]������7�0Awh���
�:g{��/�V-�?����%1~i�z!�{)ɓJ龑�c�b����
���r���D�֢�k�i�B�d9�L�IWD����Q��8���Q��bUvt^���6A��,���I����|�z�ؾ"�vc0�S������*�`u�Sf$�2\	�ת���������C^ZYhW���'bފ�Oؿ��~�㺋���lTƔjx�<�)�	�������Py5�R+����k|�ح�����T��ViH#�?�5���X�����	./*�F�9����"H�D%O������(ꇢ��A�J��3!F#�v�f�6��6#T�����+��W�$ �`�a�S���j��a����[��YK���g�ϾʏȢ�r	P�	�-5�(���.���mVբe��̓<1���>C�I��W��H�
��0�h����g�F����Z�c��̈)�1�b8P�t��\�K"qH�.���|�u/c��xoL=�V�N��*E�I������X�a������~���#�h5��[s�����]��<��t��gg��mJ~��<���e�u2>�~S����"#E����?���:�wr�EB�։{F�&Mf��#���X��y�]3���ion�"�� U�sB!��>i�P�ަ\�ƲF�R!�n�
�B�����
�X�j�7�6e��BY�W�D	J=��ߑC����Tԃl�R�����gz��T��*A�ɷ���x��h6�S`x#�}�� ԅ�P7���(�\�n��6���}d�7C�����@�!��(�ޟ�|�fz��ç�ˣ~H)���s�w�r�Q�w|���������Ƕ�@k�";Ph�F��C唦�|O����	�q�M�RZq�zN)�����^8}A�)��z`E��!r桏?1��^)ƿ\�㮽TB�s5�>��c���tY��{	��s����9�(<���H>�L,���-�� 52;РK��*<ݡ���;�+���d.�a�C��קB�o���Ӆ8b���z��N�T�W��5��(��0f�V�:���Ꮡ�ɫ�f�>��k� ���������x��kՑ7M�3s2k�Wّ(�@A�kuT]�^���>]�aXF�L��yF���;2��}�6����F����7>�� U(w��j�2/�k��5�GS؋ά"��[��=�BXgU1��Ǟh�pܹ�%��^�32j�קa>T�k�K�����
9PI���Ys`�L	�����F��2b��� �Un��9ZW}�:���m+�1�Q�۷[�z�/�V�������d,!��B�
����L�ml:Ka�N������^�^�E�$�+�������#�ߒ�Q�\(QՐ��kL߄��t��)��/�����נ�`�^�9��r��`�L�r2�V��_�)����*N�J�A����!�`��k@�+�.�����/I<��$�r��_ۙb7����d�RV<�UoU<n,�6{+�z 7,���V����NsA���(^p��<��,�dh��z�b�e��gpO6Y�8�r��u ���J1�@���'_�=�l��V�iWZ��~Ǽ2�k��d��؁/�.!��&��Л�V�)����&�m����]�[�"���Ec
km����>ʬ�m��}Ѡ"��&).�߯�#�o�����]ݬս�Y�׹���=��̌߿��˓s�}���u;|�G�KI����7xӘr���)Q�>C�m	rI�4��@�ݸ�Hd��-�2cQ�Χf�3����%Oֻh��%����iU�\\c��ax&@Y\��&�����^j��h�z�7s=-O�.��)[t�#�f���މ�����+V�s�Vmw֗�C��Uǈ+��|t)�3u�fG�r[�q�V�)��^��Q�z�bU!_{�k�;�����c_DG�2��K�;���i��e"k��3�������8�O�K�v����tF��_`�t%uv��I7u�x�+[�Ꮅ(�0O~[Kr?�$}錿Z=�Q��$���r�F���)����̋��V���	zC����E�6'cșk_T�vE��Ⅸ�(�7e�e1=��
����#�|�B$ �nG�YIw@���{�f�� �$�Lz� ���t�%���é�B�5e
G>s�1M�j/�+��,�M�6{�4'To���6��3�P�G-1�E���u3+��OЗ/+n�R�-�f�4+��v
_���:m��͐?�����M�63%5�����N�,�Kw4|ٯ��1%1o���l�y='�f֣f(�AsV����k�㫾u�4�;PemWӡ�)[X�a)Հ�M�sT�tK�o��$�+�%���#��1�D�`��$>X�3�g���<��>=}N�	V���������<�V ���� f�Z�����CUN\�"���^�i����n_;��׋�J�J� TX�D4Z���A8�س��}���qWc �>��5���b��X9��񼏌�q��G}Kևlύb��&E�	ҭ��n]٠�}H��[-�a��/�![	K	G/���HΣ/��h�t����+E�^�´�7�D�M	�L���Þ���LA.��L<d���j���v�;$�}���2l���q���]~�HXx	)l?O�;y� l�`d�6D<��ɫ�6��cJ\�2'�z���dE���+��?|��R��7/�v۴k�P���P�>z�zZ4�2��{|}�������WK���	��i)���J��V��G;�܉9���qRj�ӛ8�]h	�Q�r`�&��)&GmϨ]�w����=���7m�;�7��R�C�:����e����=z�;wL��7�|܌g�?m�bER>G[�g���[b��<N%�S�������~�o޺�y.����O���@M�=�Ks����{,�����Pi/�o@H��&����y�q�����F�v&T���qr�����EDjaD����8NAPƎ�>�<e +�ҝR�st�wU�G~��)��8��w{�1{����AW�[�&�7�7%��e�����Ў%��	7�0t�G�;AG�'�ěx�ZE�y{Za(��d<�$0\���c.�5>+���l|7~����K����	�5���賡�L�">�`��)N�V���[�'�\�~��^?�b�j��ݞ�32��P~FN�MZ/!z��q¤��g��?uW���!�Zo{�rU��W`�B��:z��Ԝ�❭��ɼ���3�j���"��w��`��\���F��jr�`���_������k�n_���W����Y�i=]�D���lm"�4%Q"[�|��VE)�P���a�,c��YU�z��gF�Y�cl���ڗ&Ṱ2��JE`w��R0�u��Lq��v�w��E���{��;�0���Vs��l�~�|��c�c]M�.���_����;`�dTf�C#��yvI��{���Lv�I�bYqD{mv	E&ס��d,&fO��rI�qxP���*�^3�P�{�f��xN=�*�p����6��T��;2�]���ZI���`W���T'&co�ZL��wdxdO�L�*�	<Û�/qP�_��԰fER�l��Ɋ<;��r�4�ߙ��}~�uu$��??299߶�݄߭��0���.=�*f3��=��%��2�IB����lK6�Jn�[���mՎ��˄K��|.�����%��Wе[��;��c�`�3��;�<�)zY��L�՗�8�no�D�3�ȏ�g��J,~���) �.�.��rpi�^���jam�H��#�2�� L��bڅ��6W�v�H��o}��9<��kC���ק'�	��~���#��>�WU��X���u̦��Nܬ�s�l�[��p�,�bJ{!2��|&�������"i��o�A��4�����c̰)�V�)�>D����f+Wr�Wx����A��2�6�{�.JN8(�wĘ_Jqٛa+��(IǨ��_��E-����?<[�8j���w�	���hS�e�Z:6�kS�<�2�.�?��^Ig)�望"|��C3�ؗ�q�x�6�_�����~��n?��9�u�
�ҧ���5��ƆT��2�X���ݐ}���W�$Pw����b�'yR�tb����0�`�ɿ�@T��=p}���d!� ��ô��!�'��fu Bw�p�	�H�h�}��y�^*����*���V	Ɯ�c�Pʃ���cG�FC�E�k���"W�ط���fʁ���zx��A�������d-�k	6֓�6֫��� ؏�S��Q�[����G�@ѿqt0�����PPIG��M�HxK�~o�o�cX���	�^��@|j��>Z;֍��J�I4�C��2�4Tf<�I���L�07�������Ke�{��$�F��#3۽�Bq�Azq�leQ�t�W�U�I�\���@�ť�C2���H��b�#��ڟ'��-�7�w�+�dS�{Þ����=>3۶c�7l�/��nǜ���AQq��BI�$�ß$����:Q���z\�� ���&9���oW������l�8��}�P�ӭWrs�L D�����֓ܝ��N�vϵ�����s],���F�J��j\<��n jŸ��s��'�#�XJl������p���̀�͔��LtF~>�|������F��J�/�+�]��V���"{���1��&n�~��V������[�?���2���3�lz�2�@��ʕ���X�s��.�7r}l��k�!�dH�����ɫJ�$�R� �!���\�D�`]���Q:��$���n�}g��F�D*&P̟2�K��(����M��<��}��{@���� �f���9G7G�CX���ߠ��S{Q�ZY���t�d\x�k��e�~�\Q|��S$���7s!��K^��O6!��2$�
F��ì��A��w�R�D)�c7��+��j��3���'�2gp3j{�7%�
h��r����W4f|MKI+s<�C�<���|��*�U��W��2ԂFۍ���"��Bs(6�m'M�9a��n�����{����RO�s̪#�PI�R�c�'n������{��[,d��}�C���04�o����\���a�5?ro�`Z0RF]�B�L���+�D�7�#�I,l.�+�$sOd>�bv/��:�+�3d�7Ʉ�]��3�9��=evz�^���*X��s���;-{V$�L��yYҵ��/zi���P/6�J�&��!|��@",�Ҡ�:�3ӯ䨁�/��~2�@��c�ct�?6=k%��h��OEɭ-P�Cl�K�M8�w��0,����*�ɳ3T_�R��7�j���K�ޠ���%�
E#�F��G�-�S:�j�Q�����eGs���= �ŭ�Ӈ��o�꣟
>?^��+*��k�����Q��p���dނ����ޫ:�:/������4r׳�`��>���^}�g��|:<��m��_�}
zҁ^UM�-k9��P������m-Gڟ�⢒~��(���'�f�>����Z^�z����N���w;_}���������WߝU�.�S���A��3��)��5�e�_��+�*(=�����b�`��~�`A���7�O�G���al\Ϳ����E�4+	xa�q���coǈ��Fp�r?�ƒ�Ϳc$d`Fa��[Eki�M�N�{Ze�F�s�"�
��:��Z�8!I+�����T�x���_C��܅�G������H�W2S��F�-H��2�r�}MW�r��2��2�b������������Q�k��Yb�Fe� ��}�oa��>2��wM�)�@o��t����Q0p_G=����.Y��;��}�+���_%�� ,]�a1$��E�i�m�kH��]����t��4�!����������S�9�B�{�rvwԇ�u��P-r�~A��Va���$�@g�h���U�:� �U�yr�_�(_X��( aN��~ղ%�*6���@*�u�����[�-UC��l]@��"��ϰI#K�`�ShO�&�4��{(ߣ,��8�z�<Mφ����$�����Y�܏���-C��X��A)�#%E�e���4
����r̽�*��lJ0�#�n�/�����������S��GB�h�����ް4�!����hUt��k�jR#�kW�@vϦ�G :ֿ���~����o���x(�@��_�E��`��\~Q�N��h���tZ�,��BAõ�Y󖢫�������C���*�m���c�$��2��=�T��v�%�8jWj� %vL����@�/��KXn)���; �����4����o����{�yI7U*�;���Bg� ��G�\+��N��f������5�Zgl�W��9 ��6��XG�eׯ�IKw�*���lU�?g�*A�'h���7��������P�wg�/����p��]�_`lI�tf`����Y���:÷��*'X��t�R75)s�(R-<� ��Z7����S��/_�L�{+��	QW��d~�{�/�����8C�۽�UP�����B�Aݖ�}�|�Ò����0�.��n�g;�C=%���=n��|��\&�V�![J6S�������;t��+�Z�!~�װL<8L=�l�e^����o;:��i/a�_�n�#�e��F�ף�͠K̞�ݼ�����X����S�f�bDl~��%��?yj�?m��?U3��U]��(�v�_@��� �3�`�%���~|�,� ���9K���Å�K��7��29����zI�4a��;P�q�`�ڄ: b����������\��DL8;����>���/�j�M��`��gM��j�;vc��]O�%<E\���Q`����S�"%5��K"ٛ��O�oБ8*�:A�	��ǃh�q�>E4Q��+"xjI@�/rBfI{����t6`�S��V���ʧa%H��d���_4���?��p����b#��I݌� �z���~������+���_�1o�y���m���Z��C|\#s�������J��7��D�e\�u���O�;6���Z.q��!�uj�s:��n��י���JZ�H��ƴ���L0v����ܰX`B:�ro�}����r^r*xCen������Q�#H�UY�i��s���,
P!�}�l7d��Q:�������	��xN�+<�]k���C�N�?J�4t�V���/0������
�G��Fl���q謙G���z�j���md��0����9C���^����OKN�3r�}k�\*w]���A�2�+�57ݽZ�Ff|��"��*����#t��g���	�����G扁eP4�{�U��<���3�[�m�#��������o�����	��o}z<T�����njU�/��=�MA�/����Z�W+xd�d�R���;8oPJ��	^�x@��ZF�K*)��`��c�,`�G�r|_����n�]ė3��e���Wp���t
�}bj�j6��^�$f�/1���Xu�xs����(�mj߭=����|C[O4E�OH�JjЁA�|Rf7s��5F�-�R���Cw������������0Hs��Lqn�0��a8�4
v ���	@*��q�߃�!�y�CI����Ɨ4q�\ft��^1s��WܩQ6��B���t`t >�Z�ܱ;t�^e)
�߅�~?)��BX��j��&gJ�샷�[��NFp�>	x�W�l�2L~ЈzMن}@��R�"�b�� i�nF~iDN��&bRf�3������xS��c2���_�� �وS�����xb���⇬h�ٛ�BH�6��U�7+eTOhXT����� �Y����1n�w��x��=��sP���D��.L�����O���qo	��g�R��_�)����9�	W�4��C��B$Cr�]ϛé��}4���p�i3���g�-Ԏ朋1����#?���6mAȧ��������Q��ܺ��m�C䱛�O.�_3Jb�]��J��P�&�cV�%�X��0�0�֨R�;����l����� :��	�AwJ:�-	�us��?J҇*H�����	��pu�$��Ti���m��y�!�ط1a4Lq�pP�D������?�]�9��-z�ۙ�#��RC*وMz���Y��/g.���Ӭ�^$+����"��>�a�ȁBhzV=ђ0�?/��4�K���d`�8dr�j+a.2S�ǅs΋<AO�9!Jt��86]���S�`\��R�W��G�^=���F??{­K���|wW�Ap��±��������������0ɍa�vS���y�������>�*h����_�F�%zDۿ�M�
b�l���C�{�5�uk�QD, 
D�(�AA������.H��Dz�.����t"Az��)�H�V@�n�~�y<�=��~?ree�d͙9Ǹ�1�9VQQLL�n���p��`窎\�x�=K�A�7.8m��)y�6�W��߿���[t݋��tM�v��ڳS�@W^O��\�EZ6",������ �� �a`ҕ�kŀ���6N����r�8�
�ic���Kqhc.@G4 넾��]jbIR	L">�t�!�o�7W�۔^{�a��GZ�N�m�K��B�2D!�h)����*��4�!HsNE��dUZѿ������77�|�uI'+�k3X��D{Cp[A�[��m>�w�f0 h!I��@�;4!E�z)=��-#-�"%;ao(8�7���j=SD�A.!��@�uP3i\����X9��xyg��	"CV��-�Ƭn���,b�H�1��S�y���l��"�f`����&`�O-�(� y�7�p��w����݈��ZI[�r^���~��� �h8���_��aj��Ͼ}� �&+v�Z���H��IӚ�Y��P�Y���sHEj�y'M����'���@{sF�_C�?|�|����Т:!����\!����.�}���n�.dĎ��_��-�K�ۚ���$\"Qb;M��d2-$}j���o2���Ë_1���4�1e$�bB|��6� K�A��O���K�5l=җ18�22��Bd�Z絾uX�%�Vl�x����޻(&����)�-i�o�� ������kMh�_>�Fɏ�}2:~>*+�Ұ��2q�zL�"����t_����9��D�ͽ�S����ʢ�gr�n��9����5��,����O� Mͪ��
��T=F� �A�@[N��aDc=��Re ��0�$��8Q�n�����`<�RF���i��:��P2�߳��`;	�V#�ACb+���1���c��N�1k���{R��� ����rR����
�G2oF��j*�v�rϏ0���<3�������#܆b?���$x�Q�&�vR	z	�9����4D�_�*������!Kڂ�h��lB�0 ���L��L {Q!=�Q5����kP��[��ɠ
~)�V��żMCU1�h��C-���Uq�l�W͜��{s5���>�V4m�z%��d3j]˓�V>�(P�7�j�̟�,��+�u	9M^�O����c��D���E�A�K���%�i�W ��`i[�/iεo\��[d3pO����@>7��(�Z���p��'a'����lQ�yl����x����.�>�m/8%�Nϡ jߌt��f����뇗��;\ة`��}9���o��șƕ����lOX�>�tv_�_܌xQ�"�2Ac�� )*t�Xv��M�t���CgP���5��0�L�M����8���4S6����S���l�b!���rV~�A�>�����H�����7�T2����b�T�N?~�.j�
~�Z���^�8I���;}���0�.�.]�V>����8iv�M_�����uXC�k�;�Uvzz|X?T
�A�F�7���0�Ƥ�2�~�U���fJ�'V,-���57��]���Լ|4��O�^Ox]�s����Gl0�W�����'�X�z"�c�\{l4DY��=s�
�6͗��W�tw�A�F���fgr�� ޔ�����u���楙Uv�Db�lo�a>[�A�W��a ^�T�~���w��[���X�=`*'	�,Ec2��r��/�$Yn�Fv�6��uM����JX?�0:ok���j_(��2�lv�b+�p��*����#��<� ��{E���Q�o�h�Z�x���0ޠ�}�bԒ�F��XD�� �'Q$,W{ލ� ̎�� �Dl����4H���˓4}�.2��Ǯ/˝Q�H7�[r̦ͨ'\-�R���Ƣ���!�MS����0_�'���UBͤ9�N�ϊ��q������RU�37���k�e�ڴ1q�b���3�@�XJ]g)cE�:}*����2P��)&jv���x����h@��s���s��A�,�䅸�WWf��M�Vs;;b��%��tԋ�whZ��M{�uB3���d��]�` Z�^(
��e'lz'��r�-06;�{�R�-e�J�ۭD���JAX��@�ǮUeٮ��,��,r$W#��ࡧz�f�R��I˯�`8B��<ǩ	�ٚ����z:��E]X1 C*�A���Q���Q��d%���"�~�j)�͇���s<bZgfh�e`YZ��bޱE��l��B&�KI�,��m�˝�~�(�]�3�RƂ��,�fx��7x�=OOU04�<DQ8O�K�m��m�q2�Y�]��+;nv�l9_uԖ���;�U�Q��=v���j���ڻЁƷ篥?�s?�\W�Z�KY٨����6�c��OZ}�Tf)J">�M�7�7NN �B��+�:�ٜ��U~@��� d�R ��$pk�J����X��M�$2�@]��1 U6��k(�R���ʏ���n
,2o�=����D�k$_}��c��DW�b�E�����k��PҰ᥌����-�e�{%{�^����	D�����Y�Rւ�Bމ�Y�1�!0H����7�W�`���V�'�iU�+���E%�]F��(\j������]��R���Lp�pϞT:���*Q�T���ܼ��"Y��D�3��֒���?������~s�2��zBZ�0��4͕<r�m�J�B%B��g�q
�j�5T��b(��M�l��d����~h�%�Bc���}oa�Nw �s��/ �K2�nϻ�[j��VPD��x9��D�����gz]�����������!�`F��� /��9:J��dͱ֥Dqy2��.t���(�30gjG�����] ��q:a�O�1�Ϥu�Ev}l���3�y|E�ޏ4*���EHOX
]fy6�x%V�_��V����6�(6i�X�P7<|sw����U�����}��l���]ybߺ�fm�97��t�>Ǿň������^�� )E (h�돣�0E�m�#�üv2z�3�X�}�� �R��x����Ư�9�����q���쑮���Oz�ɣ	�	S
�r�b��������uxY�CQ��y�#�
����+�C�����	U%��ؼ�VQ�#.){��.�`_L?���ʕ�~Q�"���1�us���NXF���>��Q�Jz�ȥi^)U�o;�X/6��Kٟ��S�6.��
m^Pc�
a<����x���j%y����J�_�~\4"�c$��2�:Ȏ���Ӱs�dC��Ş]{���2��ݥY�o�Vg���Ê��q��*�Zǐ�l:Z�������c�|E8l���E4`z\��`�{���:f��CB������b�gUЉu���o��� ���>�D&%��Ձ=�o�B�����3� ^<��-�����I�-�8d�ez��TOO/�0��&!.�u�����=|�Kl���ټRE�WEW�T�"��e��b��-,Z��~s�KY�G�nTE�یL!?@���L��=��t��=�~#��q��>�ĸ^zn�1����M�o��ē�kt;^J���K�~z��F��˰�r��ɠ0�,O�l����i��G����N2g�̎>%&�n�$����_x�[T��~of��h�ゆ�6q{�D�uO��M��(��;X6�^���J��~��{MU��1v@������X�Z��ު�ҘqKBP˕/� xW�O9~*���OQf�)������p�d����R��S
�R�T~(i͙�WF��@��4��o�MAn^��FB���.=Ӯ�@�kʺ��fa3]����4��e��vޗ
�?�M�������}ac�a6�hߋ�엡>���&�`���_Y�u�[ �0Sޚd�/'�u�,�b�I���L� ��n�n~����r��z5աQ�v`��>���'.5���*A�
CSO��
[��u���9� /=��S��������@5ׇ&��d�k�!K���j U���\�f���Hk�f�>��ۏ<}y�Hze���W3�SQ�[��b�"���E��0ٰ=)�`��W�@ÄH��SZ�Y',Z�
�4�T'lʭ�Kg��]��Wz�f��w��P6�	��M��6˸�����S9��!����?�
�9�Nx�7��K%&��I�c���d��}0`��Z���rx qm�Z�"�38X���U�w��ta�`�}SH�û�.��m��_��q��5�d}��������K S�xy�DJ�3�w�AhΔl�8$�==�<s���ڊH3�[n�a�O{3� �� ��&���=�r��o���L��tY�|���m�𒺊�nN)L2�B��7n"L�IfE=b'�o;�Aq_$� C��q�z��&vC� W�����g��L�5.Y�O��K�,�j(xU��o(�v#Ϸr����]Ƞ3W�ש��iowc��z3��J%~)�c6NA�4P��֛�Z"kM�����J�u�J0�y�ud�X�� �kc\LY3��ss�)p�р��@�w��(7jo�h�����9m���÷n�6{�P an`>	�r�ڛ�U%���#�T�?3*Mp���zx5B'��K	@3��]=���_�"[C�D��0��ZL�B6�0Mz�~���������YȒ��� R6����+!]],�o�h;��9^�S8�}R�&��?`��C#�Dx	͏���ư�$�(B��u������z��g�.m=�Ҩ��T����ƙ�2ȫ��$�>��xE��"M#��b^����eo2�p����p�0�x:6�S��1���=�k����ňG�U�P�F��l�qЗ\L��z���zk�t��uE�t�l�)e��$�ÞH�a�N*C/�	���l�[>ED6�}�ڵl�?�hu;[�����F�D���1�-������
lq�^"<RpБ�x���2z�Ma$��X�P$w�!ߣ'�V��b����g��	�巘�xY�nU�e��E��ޤ�ݏ���%`�����-��ݮxУK�G�\9�q\�+�ܽ�}I�0�n�_4�Ǉ��"6�9Y4�����Q�C�ԫ{������_$��ī�0�c�,������9�p�)��W�y�O��V�񄆈]*�8����cA̱�]�oE�y������vɴ�]�4f�?�j��[}1�����)g��#uى�-;��)C��s;B��1|�YTC!�����?b���{�}���_r����{� Ც���'()O����eB�NAH�܈u�c}�Gܔ4z�'�p٣��%,���)���pX�'�ܑ͇be��Z�0E����z�	B�c�ى@�|���G�@�ls��*��=�*|��K�t���Gm�=:�g���Α�~E��59����p7�ϖ�=��3[�Y��ou�V^�6�/�.=�~��3)� [�>��O�a��Z~���N�t���� �s"�0;k�N����Z����@ I���x[S��m�B�RP^F�邅	�yǈ�� qK����#���e�u��Cgn�h=5�y���70��F�4w"��H2H�ė��g��� ��G�7���"Ȩ�]̜	eOOܭ>O��I2{�R����(���&U� �!p���=d�M!l��ώ�L��f`�
�D�Hu#��G�m;�~�^o�08ٮ�p�{It����:�:Z��6�a�>v4G��U���ᡫ:u�vV�lY��;E��I:���	��'���_��~���8 +��2���-# �u~
l*"�{�7� 4	�**��X�j��2�+2?aϡ�,��5z��YOO�F��gЋ�J0�S�is�8|EZ�r$�ĐA������`��W;��#?"ܢ׎�H�b�8��A��D�a4i�:�����M{�"���K��7d�蟢���
�*�Vu�^�|�����s��$�������*�m��R�\���4n�ԗG2�
{F���g���Q�"��O��&HǱj�ۥ����+,-W���+�Qc ��M����2h�r�r�_�K�i�} d�CL�9�&z>�D��;m��/K���E�y��\��E���vL�)+�X����i��Y�������U�RL�g�s�
FyCջܗ�:�Il����ɔ�m��h�U�����$M���f+�2i�~ҫgկ�ʣ
�+z��a��o�-��$��.ֳ���h�Q�o�L�s�
�ms������\5\D����ABNs��3]�J�9�m{�ٮ��v]�;;5
�=��_ë�t{ ��z��-z�C.���p�7թ���1��:���8mHY������K1\Mӣ�'���gz3؇ZK�
B&z��?~#qY�2����޸\�Ixk\5��)�;v{��Y��
�d��X�c��̓�AE#��l�f��a�,�Z-8��.� 5����q����e���~����S+f�b�k������Y8y�VtX��Ԧ��:�c� @c��U�8X��`��{�����At�5�Q���$���&E���&,��x^3~�����;�t���[�5E���KN�K�%���F�(�"l�E0q�:��R� ���H�	�
��=/^Ci�0G!��&�[��f��w�~�~���)r �~��u`��L5KB���gFm9�'���ɠ���@c��9n������n!��fe��q�.��'�I-��G+�٥�����*�M2�4�ב�b��"&��_4>����ސ�mŇ;��8�P�i�#)R�]��ϫ�5טb���$��j��.Q獏�ߩ��P;�J�����V�$ʯN��w�7a����) \2�=�K�)�����7{m=8�����=�D����o�>�ב{X���v��ZD}O���w�Rbc�G�s�_��JnƆ�[������t�c{o\�} _�.Q�M�".0�~��6�7 ؞ћ��r^#�n�׳�s��Ic��ۯ�2{�*��;���-;�����*٘S"�
���
K��T���K˂�� 9���I��ڝ�e�5�T�,&�[̐�ߺ�_���J��d��.|��:�|��뻑�/c�ei�دA���tf�]�b��޾<L]��x���O�zܟ*M4 �W��|Cs�o�����a-�3c����=�+.&��~[q�A�9��?"L�#U�������),[O	�ł�����>�j������mBO CC�+�����AO zf�@O�|�.�vR�PY6��C$�݂�8?V�{��b�O��ڪ��t**��}��L�p���n��{�U�I�Y�'�Nˇ��G�c15��K� �M��\�89���*�A�U`�	�X_E'��1Lsb|��BmN�7}��[�K� ����F�����Z���p�"�싉�T���,� M-[!�d��_��8��6��^efm�e�!��A��ͱ�T��ʪꇛ�4Թ�=O+9��*���-�uBn���:'����7�m��E7�ǯ��+��0���)HB����Uڛ�1�T�շX�Md��-�)�خ̋�飳u�$)�²��a��>*)���x�C��JU�v��6F{Dx]3F<R�����9���Aw*��b�
f�^�놗D�fIJYJ#������:�aK����+O���KAk��V��nI*ܵ�ԵFÃ'�����`;�S��#v�J_�ҁ�<cu�Lx"7iZ !�|��$D(��]u!�7��W�DY?%�b���i*0��7�,������=o`�.̓*}INf杔�A&�H����U&O�ҫ�5��No�O ps�&`� Z�҇�[��/����=<��pn�_�*�ؖG1�#z:�.�L�7I"�F`Bu�v+�ٻi��N��C5�����N����	1�`2�q�8����[�y�-�u7�	u�y�/�C�A�L �w_��ٗUF% ���:�;e���ձ/�P����I��[�h�Y�Y�����h����dSq�����C����8^��C:�疒.�>���DJ��9B��Xn���s���VߪrZܑ>Wֹ�J��@�]r�;�1=A�qf�\�~�F�2_||"&V��(��&��q�E�&#r�R �J4��0�'���=���o�ٮư:w�fP�,� _��36�8��!w���Mo�l�j��H�>�����t��y�&�k���0���Q}�/�Bt��:�d�R�,	����gpOPb&�_l��1��}�	M}F#|���� k!dPWh��hK�Aj�!#�q��h{�CR˷I*�'a,�	�N%�n]AM<}�~�@ܒ�s#�c���*}�k�Z���Aa�Y�Y5>�ă�`G�����?�^-WKE�*��*^W=�V�d�9GD�.�:��ມc������,��&_w�˧�[Y�m%��}U!��:�j(�[}`��U��H�y��8x�V�mR��nNV_hm�;aGk��g�y������V6�]�U�9-��նf���i�"���m�����"WT%)!M�%�||��ׁ�K��~��E$���6���קw���|�@;%[�����4bց���h����I�J���\��Mψ7��h�H��Sl����5Ulo�.L�Y�^
Y-��� �=fS�M��lu���?-Ct���'v_V)�k��̥�FWs?|��x�5�k��7�d�u1��i��U멪��Q���M�?�3��3�-�)*T#�S�be��-����+��p�/���e3��s�P�	��k-i���D�o�u�hf{̀z�IEY%�6�2�`4��x��P�p]�
_��9vR�nظ�U�h�	�_��6?���H�?R��8��1a^��A��T���A���~�PJ\���&���8�D�o��C>ba�z�ؙx�t4s�n�����+;��7<w	����gw�]��K���j��?��ڰ�dCP;��ӡ��k@k�*&r����>�((��B����oR_*)?��gc<���{�j\��B����v%*�lg�[���JuJ����z�/
]O\0I�1���4�� �\�n����2s�4fb�0�N�3���7IV���% O��N��A~�껑���j���|�y��4��LW���LW���� �e����L�*�E�I��MpQ��P�C;P� N�%:x*�דAN0<=�&gf=��h(:\~q��_�u���^��7�'���#q�9-�J���i�9 4�<[7[��|�k�����R���ܔ������-#��f�.��r��P�+����cc�|�f�5�ͩo���;�߷5�EԜ	�a��:�/aʯ��=�yI�V��}�����Ԕ��p��AD��8qF�����1{����,^T��F��I�V����V�/�o��/h ��-)̔>>��V�G��c�?�N�;y�<+-w@�e�w�5~AYU �4x��A�]��B�25�Gp�GT�����Jp���{���}G�y�{�#?ܞh�!��O c��uyA�+(ד�o��lV<Z��J�(yC�v*
�z��}��ױ8盾a�nb���Bc/̙C�"p�wx�,�}��J�j��O���9�*۠�S_�jN�_H�sR%P�x'�xO���#=�i+f	��)G��2���֘��j��"��څo��L1����~	59dЭ6717f�Z���	Ǘ�|�>�[y} ���%���FI�l�I���J�w�N	\���Jm8��,�k= �ZD����9ii��m2���xp]���N����LP��J���*5�:킧IP���b���Ik����k�",��sW�ֱ��:��(��7W����7��Wp�Y���_�A���c��]�v)m���e^�ABn1oEn&�D�����}y1r��♫b_(O���M+sk�D�Y2�3��L�o�@�����>{y������;�2p�zw�2d�A�x����n�g���EGZ�<3NJ�����Ƞ:Y�J���"W|�o��k{-���\��Ӷ�\Z��_s����̼[���(+Z������_)YY���;P�F\�*5r
�TF�	�=t^Z����˲`�)��S'�EgD֞Ek׋�m�����ArcG�>"��[�t� /��V�pm�����S�U���P�}���J���c2�Nǚ4k��`$O���b�0����R2ɦ�4h�̶�K����[q��3��(`�� �<�'�P�÷74I�-���~�Rʳ�d_7����3���'-�b����Ns�����ޥN����^�M9�V||�'EҒ�VFI��p�n�H��-�t�R2��HכHq��t)�~mvH��ȱн�����%����븥������gO�;}��jN�;�_t��5G#��`���@a�کN��.�}4�a�$���'�����Z���o�y*�WNm�9[�{���I�^�5��U�vG1B�d�4ά�A���u5xR��@�\J���0��,Ϝ���.�Q�}��\*��E�4r쉸��/��f��dt,l�1�݇�P��!�?����?e��2���Y�y7g0\cMz���<[-ʗ}��gVo��v���pMڻ�`p�����\+�b*���u����u`.ss�S��tҝ��[c�.L�A��Z�ܵ��Q����,j�<�
׭�F+܆ѫ�Qɵ=�wcz�7X,x��'���n��5"�d9��@_�`Fe� S�(�g3�ہɻ�-*!2(�Ȗ70�zT����Cn?�[��+&|�K=�˷zxfQ�j�[�a ����U���~��r�{CY��suS����ߜ��, !�=�)~�1�n�rg�;��8��]�3�i`�o.��Q��p�5����h҆�*[k����CdPA���c�]؄�J>)KA+�̞ź��ɠ��/�Fw7�13t�=,y�f��T�$}D_ZP@��B��V���YY�f�`�l�#�k���x�V-܍��������]C��.�δ$��v�?tob]��"��D��I��f�nP����:����(��o���2#�EeRʫ��]��K2�.p�6�L�A�tW�)����w��w>�Zѡ��ҟ_j�� �	�!�k��Y���� f+�%Em4��C\edꢓE�X}܋����]|f����b���=��T������ۚȸҐׯ�h*�إ";߭����_{����N&��������ܟ��>��O��U��A�P2�����O�NQ2;�õ�/{�N�*��ۢY|pr�|���otT'��x�e]vJ��p]%��XC�L�Gc���3l6�ߝ��j����Q�V����ʸ��{a�u�#u�ɹɻU��J���nάa�@E+~i��*x�ܖ́Fg떃���߹�x�/�)E�E������> �)$����d��d-�v.FH�A5�]]�N��!	�DE�|t�����z�@�Df5]�d���Ի@�$�%����곃�c��ʮ,ˏK[e�]D��GM"85�^d���4��y�����%Q����� �fcy�D�MS<5�j�����+��LZL����DQʬ�gf~���x�`�4���� �g4��p���6�<
�6V�gg ���*�ƈ�>}�$�2#�!9Oܱ="�C'k�:A�)����E�%���u��n��A���D���6��ظ�A���ʈ�yaY��iy�j��7X/^���\�y�`�|K���i��<�:o�dl5�L}�Pw��<u2��h��a�*����Ɇ�7
DU���V�)ʠ�Xb3*��i�	;�|;��E�����3���1��K�I(�c���&`��ɠ�=��-0��So��P��'���>:��?�`��^ڞO���N�{����	��"�����`�r���/1��g��AC���O�A��8c8[���G���	 PcK�v"�$E	���G���_-0�:n`1��j5Gd��G`n�����2Ӛo�\6Q�b�~J҉�`�ÑA24�����E��S5e�Z�'ӹMQU��ׂ6#�C�\8�7��4o��-*�0Z��r�^�u9)��6p��|:�:�l]M�;8T�.f��/[����m��z�������������{�<M�˘J_��γ��K-���Cm��1�*D)��iwfR�K��"����lz�Q�T��L�oDW�o�O����i8ƐբL�vUc&��.�cL*՞�h=ϓ&���j�}����̕75�K��?����g ���Q���M��4Kk�I%��Y-�(���I��d*� �K��X����PK.D����CGW�Pm��yy�k��)�s+oW=��6�ZI(��>OxӦY]������g�<Ͷ�]U������0��GX.�_�2̈́
���7J�5�k���9�ʃ$9\��b6�1�7*�
��P��#�D�OI�2��kD�3� 6FD	���C�A���ݕ�0�nR�@�=��&�Fj)p0 o��Fߔ�f��<�pP�;��U���x��AV$\>��=�-�	K��y�>�i�ƛ��Q3o���e�k��'̒A�����J{��$��;>��(�t��gB`�9��Q�x���t�;�O:��l$Vn2���K�"O@6��fr"ԷB� �h;3�g����ǿΪ?sV���c��wW+ź���M��/^���G�X����hA�ba{���Dj|l��]����#X�l�.v����
��o*k���+�b���\�[Y�T��Ѱ��Tl���	ݜ�n>�9s�"�n���O�|�v �p޸����c?�N����ق��]XjqSuY��Ge���Z��'7�N�b}T}^1�f@�dZ�*���	s�w����/4P��~�J�h�-"rf|iSZ�๚�_��I�^��8��r#N((�����SP%C�(#%�7�$�	����T�Yс��VNi�$1>4�����w�yyJ]�2f��ٞ�՟��*�`�-Va���;��U��?�M��0IQ���2���a����P~���eO��һ�J/��7�=���ӬQ9�,�V 9�$�ӟ��7:Ak�$ �+F���v+��� w����ܕvq���]�$�޿�����>D�Kg6��L���sܜQ��g8�}�Im���Y��2)uW8,�,W��*��QM	0��哺t{����8������B���͸�d�3�;�).t% ���J�6�i�4��6,���V��7V�q0�[=?�Q��U�+����2�b�� ���o����Ay��>���?bwP�ăp�B<ȠGdд���B�+�"�R��5�5oJիwk�{ɠѻ��� �$b���Q�z�-у��R\�~h��!���]T�
s`i��Np#�<sH<a5H���ֈ%�$b�1��f�{�R�a���"F+%���*o���	�(G��p>�t�]Ɍ�a�xK%�����A}�$Y9�)�g�Zl��u�'=)c��1��=	�Ŗ�?��R}?��Ra��x�z�eR:O�J�lQ=Xϩ���S>\��7j�$�p��F[*�2��Q�G�
�3.�Gh�D9ǫT���yx��@��oh�	0����u��g#�.(Ѣ�0*�"Г�t�`�c���G��������nRy|$�/�|K�����K�j���tj��ȕ����l��.�?4��p�s'���3�ſ�z���(�>�"�4�<8�%x�}��`�A�!up]�D��}I�Í`�aV��[��^�:�V��.>p9�tK@L�C�S��Gu��s������;h�V+��g�^�s���k C�8���l"�c�B��@F�1CaU�3���s�,�qr4����.�\�%R��A��߽�}���ը��:$�B�麤��І���r�{��m=03ϰ5B�9�d?�t����?{��5|�xO��҇Й���8��;eI��&�ZRi��/�}6�t�B*e!��	��A�Kټ)���ЍwL,�ۉلG�; �W�SaDe�-�t�Q����{�"�6�%ڬ����R�_�u�D�})��BS��f����cা�{��qd�ͻ�����Vk2�[�-$�<�������K�,"���?�98��z�W��IO��h㞢���}���]���<���YT�Ĥ���q�0].�G� |]�juD��~aj�D�,��4���*�Jj�|��m�,ҜU��@	�aH6���M��ƅ�L�pɳ/��n{3�9}wYp�&��2��w��3�
(���ݣ�lJ�W��(�^(}�����S})�|7��.�$�AQ���s���%��7o�5��?3�O��=�t�����Y�b��1��m�xjCNq�,r�턚)v�%����u^�u���@Ǌ�mYq����>׾#��5	�]s���9O���\���q����W1O��{f�Q��e}qg���hQz��h���|�d\p��-v�};2hy�X�/�"���¾�A�^���b�Q�Rz��*�8xJ<m�S�8:���]�奁*A���Hi@�D�q����n�*�m��:�D~\!�T���S���7i�8U�#_i�{|�K�r�Ҹ#C"4�����tW]|��I�3ꪢ&M��I�I����e		J�03���;���&	m��iV���7�Y�G������Ȥǟ��!u�Z��h{A=eZ5�Uy0v!�,MB�3?�TWh�^5!�zjf�	��r<�׀ڎè�#���K9���L���s��h�9L���ѹ៓t̯��<ҥ�>���U��6dR�au-"�!�iL��� U]�w�4>�M7�<�Xɝ�~}e�VC�~��C�t�䎗���B� ?Q����ߔw�_"<�����RK��j�(i��"b��j�i��%I�s;�&F��)m��I�Jˡ�n���p1�,�rm�fxwjvƂT��&��w5��A��~�Em������YV����~�&J�`�$���lb��D-u+G�k�>�&(1���uJ��,���|�UV~1�)�7�)�1��N.Kh�����+K6������/*w�1i��4�=��GS��j��Mq������{�n<�ݠp�I���a���q�p����,ߢ��U�zn�k�'X�P"��J��b2�b':�j���ʣj'�F�V�0�~�n��j�}�����*�b�Ԣ�JH��K����I��%5>�,����Fz�*��U��N��E�\�y'��Yg�R^����P��[<k%�e�J�W����}��	v��}m.l�y[��'?3W�ۺ������G�Îi�(��n��o.��{Jh�@Iќ.o���Rc�F��%`�S��G��!zb��/z}��3!N?:UQ5� ���\Ow��e	�C/̸QYsag�l]H�R��d�iVϓ����
�*Z;��W����>,
uޞsu-~`Ǿ�}JW��w�)mξXι�Lᯢ+��an�Z$k�^�5�YH/Q��y�m�����@����_�9��~R(v�
c�_Q��D_1k�CM�*PY��.`�P �����b��)_��UUg+���پ/��8)�k�9�
����n��M߬a�O��G�r�W�}b�l��n�Q�\��X�R�5.�M�B���������̈VV���*�Vj�љ�Lw����M����m��}vu�:���`!P�Ǚ��#j%z=����:W���ǨYuf	9;����FC�;��4$Eq�geI���(0?
� ��vyHz�h�˦`�h�E<�:�,$O��d,`�?D�NU{�v���;�Oa���_q����6;r��� ~�b����d��o�S��OG���m�c�Wrx�%�5��ʗ]	����N=��{fe-��w�t�g���؂E�d�a�\V�L�ԅ�Ve!���
�|�L��nU)�/�y�Zl�ʤ���8���x�2ß�|w�0�F�×��8��� }ܖ�M@�nVe�^=X ��R;��-���%96�:��"��=�ƍy���h_�
��/�b\:V�ǩ��Æ��XJN!U��Pw�!��-R�?��w��6��ʃ�=}-F��6�j�jg��4����_4��nhJ�?�K�ȴ�뾸����Cu;H��U�>a �ڇ�PeԵ
Qڬ�;Mb�Ƣ�ۘӬ�f�u��z�MrAbF�����e�|�$]�&�~�$h�+k{e�/IXP&�<���}��W�V�/KS�q�1�?�Z� )���q=Ǐ�����q�%���ޏ�����	����{+%3����#�0D'ؔ� �P,��:n�o�D2<��=Ia3���y�N���-8]����L����']�����wİ�A�=�j��1��!}.m�3���M���Xt�?���-�&\�_SH��ȱ:��|J��F�����,�p���e�N�<����������EvL;���Y-��o��E��Gp&v"8��)��w�)�k�X�Ú�|p@��o%����0�����d*��4l�Io�v��l���|_ݣ._����|r9��2�ً�R�dw��6�U�^���͔�@��?}�����.l��N�*GQ0{L��Ǩ�'�R|y��rM0^���;�	���_j<����&����L���� ;*E� G}�s*d� i^�l,BZ�Kd�.L� 4�SE�VѤ�䌝�E��/�QD�wd�`�(Qײ�I���~%dT�՝�A��4���Ф=�. >eCmR\���T������\cL�
/��IL�� C?�Ex��
0[�����A,q�O��
�e��,`\�"���Ć8:�O.����i�&���R��&�d
zp�i�M�����9��JGo�q;s���ҩ_�Ǜ�hه�v��ʯViA� -o���;A���A�fvMM�]10��~4#)��J�(I��J ��?E�od<�­D����+��Nn?��Nw-�A$�k�[A�CpV 3/����uI��[~��~����>�?+�/^�l=��щ}c��m�dg*����R�yr_���oPp��F��:w� �ܑG�,����S��ݑ���N�����=s���9+��{Zf֒��b���\����{��z�U\��P���//��f�����GM���_���כ��ښm��*���L�b�{VZ��\!�袻�23��m�'�2,rrОԭ�&x G�}|��6�� ����J/4���6`�1`Nέ���_0r��p@��c��hc$UɓA*�:_a�JF�b��m����B�{b=�&6���l� \ɠ�����s� ��8�!.4���o�op��癎�}���� ��ϱ�Ms�8ke9�:�N�}B�y�ea֫���+opbQe��Ύ@��\=}�L>[���9��T��H����%�*����I9�d����T������֗�M�\�MΏ�x3b'4�3��%�H7wYXxY��ck���,�"�wH�*h�<K���vJ>{n��7��Eq8���yg�W��jb"�4�^P�ni�Fn�j�?�´�+���K�[�� �, 0�V�z�/�(&�Џ� mG��u<*g���'��d��8D;d��Ƹ*Q�25<�=P[���F���U8��X@q���h|#��l�k3��:ɟC[�?��<k��r�b�u���FW�_��]��9������vOK��C�t��s�i�k�u��䶭QTP!���"��tD"b@@z	��CTz�F�J�Ԉ�҃t�#E��&��K@�k��>g���u}?�L�'	ɜO��c�wS}lY'��X<��G���a�mڎ.Nd���ϕ|mH�BC�����gb�6g�ӡy�M�i@i������\%�@�i��o�nk)�����z�v���|���QC�	��z�h�� �M4/Zw8Q<��ωEry^wj7�#�G��7g<�kgBW�|�rMė~Gܑ��O��;ώ��$��ڧ$����'Ԧ]��Ի3��v�_�B�|_.ofq�N����9]���}�'.�+i]��ލ$���e��(_C�� �{ F�\E��,��E��u��0�%�wEv>ZkY�̨�y�2� /z�	�Y�x}���(�T��;��mU)���RSQ�M��ė��`�S8�5����"����h��m9��AS�?���q��ե�e&$5py��o{؟V��;4*��{�gft�yQb�C�����]��
��·�����W,�wgҋcǽtHFa���<ڻD
�����<�1DS}&�Ftkќ]Ր�8�t��o�6��	�Ѯ����T�=p�1>�jn�ĳ3������׭��x1�$����d���7b�إ'�`vر��H��|;��A�!6D�?=DMSb��gBy�b2�Hsr#x*�	;b	��D���LJ$wt��* }qĒtP�rv������ Yͱ�N�Mռ���B��]K�f�\���o���~��b�����٢H�Ⲉ6�ee�9;�GR��̒��ׁ-ȏ�5+e1��m������.�Ex�;�M$<@g@�e{ 'x ��;�-f������:KƑ���#�w£��"㾖�it��t}֬Tɱ>}�����ڔ��"���~l���8$>Q�,��g�5��n\�֓Qtx/���ą�Jk�Q=?U�&�\ߌ�U/+{⍗Y�uy?>���vY5�fv�Q�uƕR�[��ɡ�@KjK|L��<�	���X�b�9���
2# D�X����Q-<���a�~����N�����9���=�h�os��$'n���39�IwZN�C�9E��=m�����4r�& �{�z�I�zߘ3�]}TI%?��~�
�ՒC��9�~];meҤ7=��0v�+�n�}R_�!.hgϚME�X9ѥ�=��qf��E�#:8��p��Mr��:pK�L}/��Fȑ�tj!�oʾ�����S�/�ëM��ɴ`J�g)ß����Y��u�b`5�KD_E4��L��N`%ӌ�1�;4<�Ϸ�NJ{@�Ռm�D<'£;��	�8���x��1,�ʃ'�m�bA�����Ȓ����it���N� dq~�f@�Lw��S��� M­��0dYH��1!�ѯ�KM�y�[�]Y�5�ϋ�"�Q�I2]#����|A�h�O��?�`��c��Nn����$���K}��Qg�+}��:��s��h8�bD�Q>[|�a��q��	���8f��`[���
���:T<��jĺw�Nj��W���~����*���B^$����_��h��˥V�����/���6I�����l�P�C���]J֪�r�U3�C���J��\4X$�I#e�!���LD�,h��3v*�g�����ºU��6���D��p�$-�+	(�үܒ��l�>��J�;���AX���O�f�	�2��.pL���.��f�F�<c?�*��瑴;`?[�0��l@�Ij�.3D�����*�bM����A��4���p��T��e^*����o��ԫV��.}]�QڷJ��(A���Fռ"��Ё�h�*3�$��|����G�.u,G��Mvᬿ�Vw�=��v�=@��Vx%�5Ne�0��p�2P�ƶ�g��;��)	�.�9�E��v�/gJ.��L�.���Ý���eM����5
��~�)���өoO����tK��mY
$�C�� �f#�l�}���`��M8`�g}��FC�1Z�<�d�P�m�i9n�ģ�!>N����z�y0�h⩶�D/���r1�۱���s]d|�@>�f:Y�bd<��t#������hit���mF�{�'GGw�Ш(m������ma���/�V��p���ˋ�;[��S���n�i��f���r�Ԏ�ſRn�%-�ѥ��-��¶�֪p��M�ɾ��I�3w�+�TH�~b-w�԰Z��X��i�%�W4������������u���ghE!}�]��UV��b�L$>�o��7�ii��6����y)�������Y#[,E����ws�5�+�v�냈D�1��,�)�v�BXN�CuuPH����a�C���h�� ʢ	��s�Yq+"��4M|8����Ҳ���`����L$qȋ♋��R����'�h��}A3>�&~i��y@{�1���Qς��Y��A����l��^<�+������4~��"]�
9����po}�b�k��w2����b��v,}���N~�+VG9�3{���s�l�Yܴ��Cd�;��U���Q���y�X�3E��✖È��1�L%�Ę&и�"�wy��)zZo��_���KV=f�Kߧ?�Bv�9N\���1�
LW�%�	ۚ�~��1{T�A���Rw'5p��:yՋ�M;n|�y�]S7nv���"X�m��;��BN:��d�����};�"�Ҧ��29e&'�jJ�3�S�t��-�d�d#tp
��'\�
R��zl4,_yT�O�0�,�������9�$��X5bE��i/��̓�$Z�T��Q���u��>�"ש�wሓ������?m�J� }�����d|�ï�<S2��</�'�7�}r�:�gr�z>�$0��O93���N(q@�"��Y�<-���z2��F�RT��Vk�:���8�wX�K�	�@��7sT\��GFϝ�'7i.8i���De7�nt�ĉ�������\�'A�$��Lܰ��?�q�og,@��u0����:y�Re@-v��WeD�<�	Fr+�J�Lic��(����C��qJX\�ic��w���z��}(�C'�ܚ�Q�9ܖ�cn���X�dͻT��=��X9�&�[�]T%���fM���vt��ժ��k�Q����V�9��C��wnM`�0��^0ؕ�)����r |��*A�|��LVPU�\[�*�ى^2yH���I�&�(���a�*6�6	ֲi��i]�e�{���]q�do�R����|��
пt���P���Bݮ։��䝽+�跨��ӭ>(�%\ע��_jO}��)��7����������'�=>"N�7��>��K���RA�KqV �7Ȼ�@��e%�9��@ۼS��,$7g�-(�_{��H�a��p��b�ɋ�3�#FkZ�3
�UF�v�/� ��_�,Sj�9Ý��F#����3`^��T���/뫞�
;����k���h�}��0'��������������mk���	>�<"�N:�]�˒�.���%��G0b�~���;(�����>b/� ���Ř���%wg�P'��_��:Ǟ��%�J��%dڝ����/Fe�At:�|j���y�m�3F���"�g�~w*��/�%�bMw?[
�3]=�K���1JJ�LÜ�M��<t|��Ӌn��Z�]*�k� GZ���cX���Kq[�e�栄M��c[ĲZ�潬i�*�0g6.<B��#-��jWq_}"uMډ[Fn�Yct�{��q������1��ٽK�o2�k�nx�H��� ��� ,�Ǝ�Ⰳ�����!鿜.�d@b��� ��|�� ��Ƣ�b������Ǳ��t��*�[ͻ���vg�g�Hg�դ)"M�;�Q�����l�������[�'�	��Vdפ����^Su ��n�tD|��p'��5=���9ɵ*/Ú�Z�8a̰!���}��ѹ��|vl��-�N2��>��.�ǐ�w*���Z�}Iŵ��őS���0��/U�C������Y9�������۰�m��H-\%A���ȸ���p�Xaa�j\߃'��:��*�.u���p��I��J�W(�C=��+*F:	�@�/� ��+����7�3��������sp2 �  @B}������y\�>��QL�
�|�f�Iu�����o\[��{���dv7����>0�CPlu���J!3j��x�I����,��������:�>U��}��%ـdJ0���y�T�-ڏ�k��/�e�"�=�5�X�S�$>�ڹ ;D9��sv�t'��E�6���HZ6Z�.�zq�5U��x7�-���&������"�_o�����rv�T��@�Q�u�}�CR��$A;Ӑkc[���G>�U�<�syrѲ_R-�}���h����o"��_D`2OFNF0�KKTJ������ݨ.����� 5�d��v��S������0a֎��M;x��ܸ��	RT��c��2��H%�	BŚ}���mj�� O�x@x���qW{K7��`�2������a�,��d7��GN���n�c�nsa��Ǥ�wK����E�_�6t5c&�S]b�\���2�<o���ki`w"�B�tl�8KS����Xc-\�2b˳��j�m��":�ICZ���a#�q��-��%�D�P9��D�[O^-W�zt׎rg�_�������mb�D r�B1��K7y�:=�iH�Sѡ�&��Z�`&���`~�Is�ix�4<����xoi�Eio/�~��䄳�ƹ����[Ć�v��7J����������JT~�86*�s�J�b�$�)C�@j3��I����l���0��Ȕ~0E�u������>��.���Z�Ƽ�ߠ
�I��*Au�A�Jk1��۱o���l�(r�N��O��d� 0c�[�/�6n�:e���ay޸ ���z�ǥ%�0�>���E�?�K[��0��];�e��-u�R�К�CAug�,�}n��NF��ֲ�Ň����+޺ �0�����'b�o�Э4x-|wB�R�:��o�vY习���QB����ݥ� �_���XT$�Jwn�X�z
4W��������ƣ�/��-�?.�5�e��BsG��JXW5�u�U?�_�DNo'����N����>�$4_hΎ�H����<���?	�s"�����	��9H� ��uk�o�V8o�Pnj��ژkTVGq��������S�G���V��eOG�=D.���`+ ��B�7�ңy���vio�������!X�V�
�SOB�/F 6�`�ޗ}
o����p���q�7����$l�[��w��v�C�����mܱ�da��+���=T|sf���_���S��x��H�%$t6�;eꖓLZtz���Kg�&�M&����~�h�2Gy�MwQ�
���E�2�{t�)�52p��	�u�����=3�e���`�Zy
ԋ�,�\�\ڥ_�#�zy��b�W�@[�����\���o=n��5�mK��"�纼$i��'��H�RM�����#~N܁4W���y��=�8h'��vq�w�T��_&��+��}_��rYK;��y������sF���^@�lHGZ���4�	�z�;ë6i[ٔ�\���RM�|/t��f�S�a�[ox��h����(i��	v�Gn�$�ɩy�>sqc�R�]J���.�W�7�np�{��W�Le�`��}�>���)zȂ ��f�N2��g�4�" ���zV���&�W�3I�o�oړ����dub�?
�ꯀi7�Ky��>
ݙ�_�}���?r=�d��ä?
Yp�}"~� ���4��^[�,�8�a���D}�z�b8�i�}2��<E��:���`�5���Ł�­��:u-!4,[W�H$��k�߯X�#+"�%"�AK&�&��۫x�6v�p:�x����K�R#^�w#������pc;]�; E��bBK����%b��*f2�x,h���/�E��ڲ,�&����E轰L���n�M����.*��������n����p��/,�*�������\�o]:Eͨ��A�;Y�Մ��g��z�:����h��]�ڔ����Xh)]�Cq�O�9L��n��n|H�j7�Fؚ��um�n�� DOr��äT���/aI�m~ea�@;�f��0�p�F�dPAY{��oy�Fl A��A0�E�j�ǰ[x��E�
�g;��?�� [����lo�d])D�������a�X��mgfw<B���ʛY�s/!+���J08�`���4�1L,Y��<|���Rn9�Q�c�>�=dC������~��iA�V�����]I�Y���`���E�/��:��v�����X�'���u��R�󳱱g��&�8�g;n��h�խ��AV�R/�8.����7�aA��7�$�?�ó�"��`�e��4]O�?(7���z�/�&r!��:?�]uh��zH�WH����t##�WD��S�[� �VxM��8Q�>���-��h�����|���D�C8�{/��Ů��Z�<���f-��ʻ7��X�4�"�鯅���<-O+��^|�o��K8�0Ŵ}�pj	9	��~5ˌX]Z��z?�����B��W�q�g$��Vk�9|*gwۘ�z��ka#_j��{ ��U��5z�_\<�}�+@��צ����r�
��%9�f<�*Yz�Ғ�P*s\M�4x���p��.	=�q�����Rp�cf=g�H�]�c�(�����.�7��ڀ���L�N>ඓ\���L���f&y�r"�̨��V.�s���_<vH���G�%cD�%�\k&Ek�8�<�F�7\	8qI@Ɍ��+�wb���@�f�1�z��^N����Ia�:p2c��r��񅛱��!�[���г���#��w�	_?[��[iU畟�a��9p�o;�U6���v�%�fWm��d!v$+����&qxLK1n�f� ��a���x*(7�߮|m���[~KX��PR��|-К�X�x7�NLM��3������ݰ/�O��r%6��H�D-���y-%��Z!3�M?#a����<O���ڋ���+U�9F���V���i9�~����t�8<�����Gͮ�(���۟����ϵ���R�髬�[�q9��SIK�z^:	vg,��)���j�_c�x�B�#r�\7�Ma$Җ;���G_@�`m�wo.��ht��K�'d��� ��s5��f�N�á7Y�e���_�9�4�%t��B�[7�tw�m�83��	��9z1߲�4�ˤP��;��K��DzQ#��rE��vY紐��~��������>���9̍�m����?)���u�J���V�ٹG��o��ʩCm�h��uZ��5N@�ў��"'r"�	����~��q�u׊[��%��,hcsܓ���۩)�;q�%�;g{h����d��}�Աrj�;<��;rgH�`���-��)]=:��$7G���V�2v��y�̭l�=��߀4z�8�ɨ���V>�>��j��������	�5�5� 9����C�H�h�o��13;pi����X�"���Z�*�ٻY��c�E��޶��,��}��a�A9�V�AF�Y�1�)P`V�KM��9WI���Ⱦ!�gԹ��'����'�g��@��d@^E��#����ŭ��Wk�b
� '$�h�H��]�^�d���md-'�`��EM�~�`FR����17���v���Я}�vd��9Gz��� ���Ks����s��+6�
�,P�+YR=r���nKŎ���x���ի
�T��_+v{�FFB��pI�E햓juG�)|���� 
�N;!z0���a6�q��\��"���2���0��C�_�%y9_���]gۀ+�t8=��e��w�F7R�*TK3F�� #.�6 sFP'`F�����]{S��{�߬�ӔKF���㩄��:���U��3#���R�n���\:W��z�o.�U�J�[߽�Gqҕ���G�-.�r4�Ug��T�*�V�m�"���-��: d�-9=>7���{�~�հ�h2�f�<#S2�j����i�,� ��t�{ Ӿw�?�e�~f����wPn$���*�L�g!�<��tGYC�%["$lP+\{�G��kHX]fڍ2�nuy���A����k�m��n�tjB<N[�[Y[�$�3:,�w���L����W�5zF�§hsu���կ��wMq9�O�/u�z��N�_D4�H�!��9@�,r�g{ vVĮ��Y ���1�e�~�g�9��R� ��5�݈�8z����p��<iy��/���ߦ"p�챿l�1�BWߣ�݃����ǎ"^�V`��=�ם'E���o�3g5|l]��G�*J��,�q���A�z٘h[���˸�
���<�n�ȶ�gz4�u���}uU��~��m��� �|:���;�Hs�|�*�!��FL��Ig���<�_E�ִh��,|J��f�����]W�?a��?0� � M�v��:�We<��9>��/U�����}t�����|?5��ӻq�#��1P�B����W�����az����Á�=��``��_��چ�O��Xڽm9��=Z&=Ǡ|�)�CqųZn���K~G��A&�����Vf|�i3o9ߐB�>�440�4�eg�O�F���U��=q�ā�(
�7Dm�a�����c�?Ho�s�C�}�Ɲ��%♂	�P�=Ԓ���p�v-g$]Д���L���N��V���;�W���a�k�CVz�Z��`�3(�;�w���^�`��~j's�Mu����?�����d%,�R\{��x�K�F�6> ^G����qw��Ґ�i�L���6�h��q��{0R?vk�XZ�@C��H���h���@p��� �����o�53�b��%1����D�A���-�|T;���7�.�\fn��dm1x{��g:��|���}�h)�f��������f�V������0) K�sQ�����.w130z7�G���ժ ���Y��|v�Ҭ|j�D�:�<.EhH���ĊI��E��s�a*��5�5����1sY�9<�_+�2�Y<o�i՜�p1�@B�>b�29�ol�b�������jHw�!�;L�A�����s�$�%�Y���������ښ�?�.S����������M�xy��fE:�j}nw�&Ɖ����C�w��%�҉I�>>S~|E�,���mH��dv�P2���L�;$`kʼ՗���8A�#�{LL��QpH}@[������{P@w��������X���k3��]:?�Nj�N������=�
�`Y���KU\D�b��خ��|j�+d��@f'����/�>?�U ~!�R�f���c��D/"5iO/z1�<��7��"TF�n�yOM��5��!��,��?*lchnR�Fq�*Y���[�a�J��E�7��V�'�����P����� 6<<�r�� �8��w_а�c_�a����D"l�0?��s����%}�ܚ�$���rY��4	/ܱP���ǌ���H��;��Fۙ���.Ҁ�.�s]=�(5���G�]�M���<%i�rH��������u+�!�RN&��m���{����7q�)�\�6�Y�e�!�h�&];$x�&��H�YN�Cae�;Y�6�E�3'�wض	�9j�s�U6�7-�
Ӄ��Qv!Uy)l�R��"�G3�'�IƸ1$��҂��/��2ƺ{���y0�������������r��^�Q˻�}�� 6��xo�lu'���sg5��"D4���]m�c�6Y^�ц�ȏ?���oM��ז�4�&��:A���) =P	��GO=K�=�s�!�j�5ZYM ��寛�=�dJ.WE�\">,���Xh��!��"�6׻��F�SW�yK�`��e
�o���d+��=��^��o&��7�
�27��/N�i��d7:>�|��������� jLS�*��\?�]�@.~�c����	Y��UkL�22���/�ܾ��{�4�);E��a��m���ɥ72#��϶�zǍ���YWh)Px����z�BP_��I�RT��R:	H=IJ�O?Ƚ�j���"~������S���*�����NQ�з�ʻ*�)֐�9�����
/W�J}]f(��[�ǯ���Tl���g��m�X5��i�p��dY�6�|S��H<{E��S�B�������9��Fg�@Ksx��+���j�k����;���^E̍<}J��>eb=s$���S��z^��\��V���Y��D�����,Pu�7K��q+n���&\�=�r�i��m���Q"�:�{R��W���V���N�����)�I�:T~����D;+4]����l�Wʿ�"A�lv��z�����hDRu��/=�ʜ�nx�Ք��	'�����|)q�z9?�ğ���X���ӵ8z?��k8�x�����N
88��J[y;,�kw�׉I�/m��^��9�PȂ&.2��1|*�윕aZ�����E�\G�_�cZB�� �i�f�m4"_o+��g���9i��b�� �Z�7�BX�L+}�wo5��va$h��Yy����V��jZ��3/��ݡx��3l9|���?���$��K���gL�7�+ 4�}�ǳq��/�U6a�:o���8��?D�:.L �*�M����A�8l)�K1Y���¹�K���ѩ���O�ON�3��b�F^?il��4fm�n��#:]!�н���������/-��Y��K��z+ڀQ���Fh��j2-7�U��.�5`�|�|b�.kTn� �:�A�d�U�ya��b��e�t�/�H��V��;R�pa���
X��3�d�X�5��E���Y?�y�V:�K�s�x�w���݉*�DO��^���*�T�}�m�� 5�������S=�D��t�~6>�}N#�P��	�h-/�A���ޠ�Y)�ۙRR�\��!\�ӭ��N��v�H�҇��ؔ�۟�HK���-#�&ʽs��i�f�
ex���_3��UX	K�Hhc���Q�[H�I��`�Y:�-`�;��~�lc|��/ 4b9ZmW�Xّ�i���n�T�,�4�H#;G��\�F,����^E�鍢�HS���{d"$2�����{�{ R���#���BL*�"�c*��(DM3�$Dw�&_*ё���5�:"v)�� ՝���l��<�W���є���L�jT�5�� �#�=�w[���"��7�jV#�F��/D�"�#�<D���B:�=@�*�Jg��|b����.�A.�)'��qk����ZHH���!%`����k>����JF��h}>wk,lB�g����e}Q�ʯ�������M^f���DtK�r;E~ߙ5�O�:+�-ߪ��K|>��twty�L�O��j�ä���h*�erz^����|鈊e4Oݹͱ�e���n�������;�j� ט�pZ �W�2��Ҙ��_���8NeT�а�9vEM���q�����7:���
�����S8_�z���r�ɰ\�u��*ɨ���T��ҩ�Ů�s�	}�鿸;�;2<T��-�,k�a~����*�ߕEe"� �}<w�TΗ��EN~[60�<�q���ʳJ� ���5��-�T�������QNk�+���0�a��8�:�腙P�{*
a�2��Wa(r1t��8޳"r���#��|��G=Yo���?��`�-�3ݘ�CSנ��[�4&��U�-E�m������T�a�9�唘�Y�V�O��EE�·U���P���/R�ܪgc��͢Q�6o� �ݠ��D�>n/k�g"0za���O���s�u`r������Պ��E�'����O!W��|�+nGb�^��6-P�$R�6�ڗF�ZvNwT>8η������/|���%�@��pj:��.�y��NL�/=?򻡸�Z�g�x�Q�n7ͷ�����#��	�"�D*���py���d�r�>��O�=Cj,��7�{˽sF�mc�L�ZZλk<xY�v���i8s�<EU����/U��n��wL��c)`�<ޝ�O��(w���J�ur�����)�Q�l?�ڊ�����pp�6� �>�<��HL7��pZDF8�ogk�ڻ�H��P����o!z.��9�i��H��^N큼&�i#��ަ,��2Tt�<_��,1+���s�����JT��v��� ����2D�":t�Sk�z?�p����׀��$�TI��Yr�
i��ֳ�wm�@Ss���Hf�	^K�k|��<7�l�~p�U೫�~���h��n9]���R�1dF72�Ur��ыa};��{�`�6����Mj�P�v��P�'��~�3�ϙv '�#?�4�7��@�.a+�ϸb��u�������*?_�;��E���8��0�w�bhխuh#��h�Uf�X3)�Xj�[rA�P���s�������|S
W)�����=��[gs8oF��=������n9l�]��������j�s��z�l�k/�Je��5>^��w�]3⮎y�YP|�3�*��%���P1EYb:�;�V����r��"�%{��/��"�A��vZR ��	ZP�b�[���2�WD����7���ۛG,9V{p:*��y�Q�����Ɨ��\-x�Cu�'�����C~!�9i��V5��k�|��X
$�Wu����+4#"�k&a��_F�Ehk�,�GuT��sf)�������7��j2[�����'�v���
��n���u&߄��s�����o�k�#�����%�eL$d��1��<-�ߍ���U���q��= ����CF�3���$/#duy�/�����t���������`�oʟ�D�����*��{�/���k�{��G�-�=�,lkz8QYEQe�
L~��m,�[jJ�K�����M�jVV�K���ЎN}~���?LVs��`:^�'��r:�g�o��gJ�v'?�!�ȯP�@�	v���v�a�w#!j�L�<S�oA��I9�������I��7c�N��Q[�*Lq}̒L���r��Ox�O�?"9�D�c[\�BQ�+�:by�s6��_R;��*��wU��������G*`�6��t{Q���c
�Q�o�)�|�d��'�����Tf��-*����ܙ�<� ����*�'1[�;���X�«O��ܱ�Y���Ix�Kd����
z=�'�H��6V�9��6�ߥ=�2�o;�5�嚯S��&ҧةE����d��@������cz}\�%{ Ȱ���ؠ�/�O�Z�z����"4�Y=u�^�;#`����*F���)o�kF���������ǒ�N	qd��?G|����LN��ᣡ]	���z� ]�s��$-}a#l��E3h\��}���aoF
[Q�����t��#�$�V����,��LMm��{V+R�*ԕ@����|����8P�����d�Єz}����W���W�gW�����E�y������`�x��V���S�=��:)ʉ_5��������O�y �%��Sܡ:�[�"�ԅy��>��g팂ۗ)� Ϯ���@����:P��r���9��C�z�?$����Q���}Kr�䗵�S]^ �F����yH?������o�*�tG�U�-�m<�L��¹����/WX�=8g���[m.�A�'�H�:`ΟZ��=!?�|���k�]̒��\�r��~���,z��L�q�@���iF����$�pa)�1��G?t���Az|v��m�X/S�ŗqy>uJ%ғ��gF/it8[	�;����\[98,�ټ"&��woe��Ȁ�����zoh�yk7[R�_D�e���w�a�iD=S����_*���(�O~����S~��Sf$��HWD��qR|,U��s�Nv!��(Z�gF'����Uwc?��5ŗ���+
�(�����eWW���d���5,�vχF�h.u���LQ<�x�6�ؑ<p�+��퉮�e���Z�q�k�媺��R����Tdw��[�g���x��A�����fD�_�_���S�h�����	7��AԆJ=�k����+A�9�\&�8�-2Xu.RF�5�z'Ń�b#ǆ1�+>w�	!>a����5(��a��q��.3�q��N���}����ܽ�{����z,��Z�@k��/�S����o^�R���˿#]2�?��
�s�YD<�a�h��CY:�+-h�Ԉ&�JW�)�����7�
ݸBw���z}�7-1N�:�;�_����(�<��a���¯�JO�}JOFȏ��xq_�h/m�]�p��7��)s9����t<o^��S~!���5I����pr�i[�ë�l����hk�6�����[�����Ո��{����$;ͻ�. ss��Su���c��9=y����7�[��	N��i�.ү�~��8�p@���6?�a��I�5���\`���-ʢ7����<��\���(s,X,�O�4�����J#���P���Ǡr�Y���c��������ތ:�_&�L�EH��7�~�J�K6(4��&΀t-��ti}u���:-���pT���V���1���8�r��.~P�uK>�}��B���5R�p�=� �&N�`'Z��A�I=߽��kb�o+8B껞z�@U��
h��ݼ)�O���$E!jԳ�s���y��bUy�>��<A�d���a9�)��ij�J�e8O�/����8�L���t������J��7J���'�'�	���$RF�ͲL�Á1ǟ%}�6����`�I�'���d�t_h�@��h�-z��<FLEԗS�<��S�H�Z���R_�0�pb��0e�\/��8zƼ� R��a�{��W	�y����^�''��4�!�Ğ��k�T3��Ŋ3Q�+o�O�x��8h0�Y[��h��|�=�m�s{��=�)�=�ջ�-�����y����nة�	t��6��#�'��&�" ����,��߽��Ԛ�g�tw7����N��A�wBƼ�a����/t�Sh�&ԓ���mn�c�� oLj�|�g�tNT�U��ƲoHdi<{6�og�
���]6�mR��<@����}/ aļ	���Chb�s��r��$��
u'~-�\9-j��iu�t��Y2�păT���JO��Ǉ�!����<�f��;�a@���G���pJ��(g9i����y�[\��9�xU��(	7� a'@D,'�&)� �A�}�t�'3�3��RsA��g�}>CCxn�x�~M3����J_���la+t�E'l�F��q{���= ����sX����|W����(�?��aY]�֒Q�'�{��CC����>O��T�#�QQ�"��Ug�����޴����[��{7B{G�=7O+��u2�.׾��S�(�p�O�H�ό���sv׉�Rh��G'M���d��ҝ����Rn�eu~�Bjqe�'t��]��*~�+�Y=f��d_-����A_�/̧�P�.���O�o���J�0C��J�����Qw=�ws=�WM�}t>�W����m�H~��!�'Tv��-�C�����X�m��h��ZimB�[��5H>>���~�����Z�2��JXi��.�h�Z���r�/��"o}�:��x��������+����:O�Hm9Ū|ğ7���8'�|��艖�%R-12ml@7��_m2W�e?�+�U�v�Ҭ�-�ɪ�s�=ӐW���8�$i�ޯ�BB���KzI�q"B/ޖ�W:Ǹw�\:�e��O�+�̡���֯D��N_��0m>��ڍHI���T��a7=a
�>b#�<�9xDV8��Ҥ�/h���W�q�vRj���:����~6�);x�*��n׽��li���e�y!y�%N;G}P,:#��<�Q:Z|�)�r� O��9�kX�o�U���N�֩`۔5��:M����,4&l]!!*)+�kp؂��F|#zfN("K��̅����USQ?��%�1Oԟ�X��i���3G�!^X��<:�]m#Ek�CG)�98p���ZP�{�-sT����|i��lti�a�I,���.��fU��ߗQ�>�:2Ki���(M�/S�i�������X��UK�0��M���F�%+��*�TK�U27ls'�(���(y�����"��<���{._Z�����s�Ö^�у/�lq�R�ׅ���tW0�N�5wgFVr8wЍ/�|�y��|r���cj[��h�����pl��#�s���"F���j��1����f�k��6��
\����������>�2$��)��r��tEo�̊���Z��rl��%�,��/|���k�5Hތ��5�e*��%1��7n��*rC�v�x�v�O�dz,w-�ЩA^�i�Q�c4��,�]Jʱ:�0�}�(*�eB�)D�og�^��gD�}|O<��8��n΂=��r[;H�_�/^8pӣ�^+�j-��m�0f>,wf�\�UY�������X�]��r�21�\ ,��J�1�����9�D�)��g�P�7�S!�^yJ�81�2��u�)4�w/�TB�'���?q��T�k_�)�kȯ��W�7Cyz�[�tW|�/��\B@O�2@��Y"��� Qy�ۃ�)T}WkU��B�R�^��^���`�#�Y���i^r+�ћ�G���
�d�Z5�kF�L� K�2�$�<Q����҄n}�JVg>Ӎ��4T�)32��/]0���BY5^oH	q���%��A�Ò�|eDB|�'�<����wM_�)�('�1����-+W�}(Ƞw2$����řP������$���U�O���f��7�=�8�Q��g}p?��l�=#{Ϡ��2�׺:@�/&(a�[Tȍ�$��N;@�T�e)�XGn$@������]��Ҡgf��',�����S+B���?��@����▄�j�e���CҞ�`қ��]�{�,`$����E|�ǎ[Ló𱤉�@-�n:�`o7�L�_V�7�"���K�{�_��ӿyϟ��>�Îg!�*u&��{ .�2z6�~��������~�/喝]����,^����N��!To��P��sAz�kχ-1b�ͳ���;�$rG�;ysk�®���t��@F�\#d��,驰@+<(�u����y\��uW�[{��y��l�g�c������0HI�����^�)�L4sV�	R`z)�}�Jc�;���x�ÆӚ�����m���9Մ�i� ��9*��7���d���/h,Ӵ����XJ��MA�hU^��ml����K�*B1���;w5��\.)��x�yƭ���I(��f?>;�Ni����<�qr`�
�|㽦��b��)v���>���Z2���FÎ��'���b�� ٮW�;��.��l��6���9XÉ��K���OP�9��GT�V+��6��qŎ��Hɘ��G��/�S_x�U��\����\��� 4tP
�n�.D���řh׳��[V�ش)��3�S���{i[Ϟ�!�@����;I��\odu���Z�&�_b�5s�W�+�� �Y8�rcҰ���w�(�٣��E�T��,r� �����ؤ����{�5��k��� ���R"M@�X   -H��H�H�N$�(R�K�H��ޥz�HoI�� ��v��9����y��t�9��+���7)�YS�X�@��7p����a�����5񕬾���4W���?�d�:P�����y����?(n��%w�u�(�R��
w�dk/��[�<l�� ��,��F|�Mh�ҳ�V�K�����J��_X��l����5��^�]bf�+�#r��c���t-�8�;�s^�ɳ�28M��Nm��:��2?�.�1���'��_��֫<��'������_tSd��ۈ�Ӌ~<u�q�.�/�W:'C�/���4쵰Vq"�7=�������[l냛�pHj0��]��5���}_���,�~4X��(�=Tָ�#[ZO	`'�\��y��]���.��!}�%��I���"����A�T�|0L�D�C���>	n	��b�yP��Yy�^'7j3��;F(i%���(��=g7���O���O,��S<i8c����d�y��5�@{�s*�7h/b|��]�\N�$7�^:��"�6��m�{40�-��I�a��Ė�0D��	ȑ{&��Q&��N��lS���F1�ˬ�<�}AO%CE�1��?����KM�x�?[wag?��y���7�e����R�#Y��@�/ڷ+š�+űy��,�铴�#�J���I�ӊ?��������c2T�^z��7����J�z ��^O"��8�o���W7ٔ2x���^G�]��с�5�����7��M�PS��6h��τ��B�n�	I1�1��^�^��۠�*�߾�k_��qY������ �D��*���'�¯�lN ]�+��df�"�������L%�[ZaV�.p';&N�Qtqc�6.1ߏr^ �a'7�L�0Zҟ><}���(J��["Z+v��1�9���G��@]>W��*���{�?� �T$5bSX{�P9ඥn��q�%�f��@Ӑ��Gv�����{�|\���8�d�A����8���;d�������Y���M�j#����ɱ�LR�l�r�x�� �ju�/��3��ba�Z��P�-'�ٲ]�������A	��o�<�鼶A��g:��xQZPKT��fi'����0��iE���ԩﱞ�H�u3/7g��w6�l<��;�%Ꟶ�ͧ�}TQ�m�q��:/�C7
[=���������r�����S��"��������-74EQ6�6g��{�)���h�9���x˞7$^,
.~�u�ҳ��c��V�bP��zo� �vQ(��Ҽʫ�z����3�����j)/�R6�%��x�_,u���������l�W�%|en}�a�{�Q��>� B�&���(�:y��Ҽ����m��qf��'%[��h��(0�t��ٜb�p�0Z3��y�Yo�5wJS�&��8xo�k��������,�_�)�\8b/�����MA���xU]"{�a[�`~~��'k��{�ek�/ԣ��n�أ�}�p����*7�@$l���mVNd�[���G�	<[}��m��A��'N&zr�]��^�N!S���u�J��6������|g]���(�6�U�L\U�V͢h�c�|��a������k�br�qͣ�� ������r����s�6��B��˗q��
�3X�N��<�l�kݱ=E�cxّN��Wm=�!!�V�����S@�����:�A��E�SY��aåP�ϖ4����w>�����>�T�f�VaNJQ7hx�K�޸[��ӧ˔X� ��ϰ3�;�߆����mPa;����k�{�i�sj�<��Z5���%�T�K� Axch�;�X�@���,��<�"V�;�[���a�$1Q9�85�B£י�0�"��Esj�ݕ��p���9aK:�݂�\�"�5 �ؐx:�щN�/�y�F�m�aE�m4I��պ4�[�=����}��"�G�"#U�x9a8p*���S���l;����|O袁�倃��m���
����1�[���ބg,v�机�Xt.���{?��q�e%�ߐ���%�q`���.����J�W��U������%���-�.6A��e����|L����E�S<�,8t�oM�O��@ZK�8���1�6t$�<Q�~�1z�xT?K:LSK�Ƞ}5u9y��u˟��ZW���ͫ���i��Zׂ�<�&��~���T�J�IG�H��|`O��T�����,���`Y��U.��4G]��V�ޢ����e5Q�L!�A��f�������t0��c4��XyD��in�JkM'V��T�����U5��nR�>
i:�ɯe_8�q5!(�K6����a���t��ٳ)�Vb���6�#�%����͘�����:�wG�:P������ZMv�Ɵހ�tz�fXM��#�b��8�u٬�Z�������.�-���8T���m�dwbG|�JZK�Yu�#��7�?e�� �'L@�.���v$2�%�}�
Wp�}z�k�f�L�+A2H�����w"�MdI��&�&�4�I���#Se)F�ɴ��u�+��|�c��������*��"�אG�m�l���N�<V�tADx�'���.�e����̒4��ˎ�j�V���1W[KXg9�sOZ�ӎ"[3I�F!�G�-�~�������J�:2O|3?K(�~��]�F/�:��x���� o-3�TH��t�-H���{<�B=�ŷ��ӏ��ѳ�+�:l`ڵw}�Aa�e�f��|f}����Nx�)H`zf1O"��eZ��`�ß�!�h����T�~��h���i�}��ve`��֗b�&F}��Kv�W1��L�Z,���S�������׶A��0���^]�+�9z]�:�;��.�����[i����龑�p�X�D^Y�a��N���s�z,g{��*b^�j �77).&�g�XUztƄ+�n��@���"����iR!� ���҈��kq1(�鵿/��q0(ߠ�	@q������rl�RU���s1u�=/�)�W�P�w����	j`�|+��.$��?�]VQ�J�K��E����?���6��;��Y�8�+��m� D���TZ���M� f+2ӱ��<�!Ӭ��fO#�i��g�Ѭ�:�� ���'4h9�.[��$r%d_U^,��%3>��Z���XNƎ��Ⱥ�7�b�Tfw��cߖ�l�6(
�@g�VM��ν���M��u��f�y���,��(���5o�����X�����6�@$/�~�8�HW�Q,�I�B4'cp��5�m�k�,�(V�����f�������t�|�U���zF����m��j��e�����{p����/�nܻL�<��Wobǰ��S@L�H�w}��ݿe��Ԗ�����]�����x̑�J~��G�4 ��?�����MՖ��r�Uߔ�TJ�a�w�-L'BN���٨�U?(�N�eZ�b0�ʻt�7;�q�ek�����h��h��ݢ^��ΧQ�K�il�1���7}]r�I��y��{Y����u�+�� v�7�q���+u�bn�#w�����Ax����}���n!����O���"�!u�Q��&߄��GC��b��~�ub�>v���]ٷA�f
��6�5�;��p[d%���F�pku)����k����l��꭯�r,)'wHҘ���N�_i��*c-�@5�O�[eG� y�26�΅6��Ca���o�7 �?�7��x����j���eÕf�/t�c�A<>��u�_���m�HV@�5�04[*u��58�(�!9͠���!��������b����BA;.a�.�K��ܛ�����+���ׄ�����{�=^�q3��A����*?�8i��~���W���叺ش3�n����˲���"��,�eڗ�f|3���L��hFN~-�B�d �(��Y_�w���^(i�,���L�]��������\r��&��2$>k`/�Ѡ���ѩ��5�w�mAx� ���I<��ni�kJ�@��ۀ	+�#�fE��ڽڂvC?�/�'f�p�
��f��aq���?�9؁�#;�Ao���`���x]*��l5�:��ަ�o��:��Uh�a?�˿&���&&}m�w��li�E��W{��X\=�Ȫ��&��3O��q��,���Ll�hq�#��!g�(p�Z�C�A�:8:l�^;�<���~w&��7D�F�:�`�����}���������@����U͍j�.=�C)/'�y�WV��w�ʝ�a|��x螝�Ɖ%#�Tv�Sz���)[���纰Wn����+?^�/�e��l	�l������aˢ�?� ��X����@�o��%��L��_U�LC�*S�Ʈ�'�����vt��cÊd�A��m�^,�f�I�����a �0�ݷ?&u����:��ہp���ī鿣�$���ȐHhV�bOJk+l2��A���[�!/f�!W��
�Ve�������?�x�;�ԁK�Rw(�}_�>4K��&"����9P���)��Aq}�����wv6&�!P�A���̭����8=ʭ��x��Ê���$��4�}��� ͜t��YM�m�a
���>���"0_��z8x8zUcv�]��.Y2*�'w	8%����9�;{w� �K�����$�=�����6s7�4�4l|2��uj�ˏ�2��e�|�+��#$���#Jܪ��{U��RCI\�R��?(Lod⭅�ʧ��{_S�}�+��:��5���D��J��1ӓ�]=�ļ*{Qo[M[?y�S<��b��~��1��M�>���lbfj��B�� ���mE����'�¼K���������$���@�g��H�(�c��3&��|�TCK	�dތ��"���'u��4'��ݭ�3O�#�^CGg��6S#���yԫ�������u�Y�%NK\ke�Um�_�a��8Ǹ���6��iu�"���L�*I)c��Էd�mЗ1'ꨕ%2U8`h�0�
�v�xGN�ޛ�č�˱�J���2Ď dsڽK�ы����o�-���Y*���wpT���xt�w��ר>Q���!,��q����^���(�1N�i!-�<�ۼ����R��zN3���S�K����	��"��FZ�嘳A��Ҟc�*���g��^�V��H���ǟZfNኌT����2�Ã�=@8�;@VC��) �z�^�X���@GjH�����I1O�\~��j'��q09�UH&����WLh�+���f�ik���!N*��h�8�(�5+*p0<�Qaպ)�\Y΄��ퟎ#��YjG不��p�Uqr���Tn�=̐nG�O�2rz�A�P�K��of�a��������F��uS 7*h#3v&%3��������I7�gא��u��n#RZĵrb�쳐���c>���a�wQ�od�[p�3�ثC�N��b��-aP�\��|�L.#P�\�X��@��,<\S��Q��.� ��FĒp'���	,p~�B�,��HL���mv��ۉ���4�[��U�(��(W�F�EbɉK�����tH�\��_hǇ���(n+�ܛ��J�LU[<�3lS�z�I~Zp��H���kI���y�eÎ=��ӌ�@�����1<�#�����q߯��?B���9 �`�ud��y�P\ږ~jü�1F�����c7�7t\����$b꜉�t� ��-�C�t� �f����������3��T� 8*���
"x�[{ܐ%j���U��/C`�>]�-?X�h/�od�)\P\5U6u�M���WF����t�{5��--��
��N��7@�����`�sdڴ[%8���xE�M?@2��^[����R�-ѓ�(�I�3�p�å��<�A?DX��� ���Ԟ�y�v��>;�|��ߪ2�!G�~��9ܤ"�����o�0p�x�H��5�t	�s~�6yc�~�i=R�7p�&�z���Z�*��þC_�ޥ[.̑Y�UL��%jν�ԳO��͛�,�kX}q<�kQ/Ż��;F~h�׵�몔�˖��B��tgq����yIȜ�c��;�w���*6��h{ۤI�L8�^�gXe��o����EU.�u�x���ʦKU�u��ُ�\_ŗ��Y�v��z6����b$�j�.�	X�5�'���Y�1�^�+���aw��c��bҲ��,\�f�\��F�a�~=D�&��z�*�*���b�s607<?��ϥ�+2ދm��=�CA���>�4����j7���O��	��$D��,�,v�HƩ��i���ݬ:�~jT�|�)=�V^��3V�;*!���!� /�������/k3�a��#l�Ӻ�͝�g��Z�FҎ�P��j��y�Z�vT���4kP����E>z�p�׏髇Fa1Y9�'R��j��^�k�j�탗��!:�W���2�z�\A��%�B���#qr��X�`��+�+�V]�\Y�+s��x�X���g���:�t�:��t�{�"!{�8!� q�(�_~U�S��rHk\fS�`h7>�����.<��&�U)f>A��)G�b�Hۍ�ݔ�L��[���e%�1cP�s:ړ��%�v]Є�����5��Xr_0��9�q��L������K*F�1*N�!�4���S��3(�j���<�y���1�h0�veNG�J��E��֬_�`�G/�3�
S?��T�jѬx�x9Lۂ��	!�?EvIA��:c�K������_%���Pi���>"o	f��3Ɲ���{V�	�z>h2HM���r���7��٩ΓV�|�͂�V>&#�����+�'~�B���N�m�b�]��D��e,��u�詈�O"��1V�r�2R��EO ���H�DP"�� ga�������u3�wQ��;[5s��p���H�o���O]���>$�Qg��ֽz�@��z6�|p������W����p��·}���E^�s���� �6�UѭO�c������ƺq��;����G��v��-�뢕ߛ�Vm
�@�Jz�^��o��޵��_5�>���c��Jf#z�1�_�����E�q�9_kn�}��Ծ�U�\x"V$EFP� jc��_���=����#�ȅi0�;r̤:[�czH�� �/�����e��R�P�n���e͝��\�&K��@a��#@(�:�+������a� �W�s����gJ�l\�;��a�+��R&~˷�|ޣ���E�§��(�K���T�LŅ��rP��Z����6""m6��Ik��_~�m�F��Jm_PdE&���X����J����9g�Q�D��XlOY^�͘�bSf�{�Kǀ�M{>-��@�_C��B����t�!�5:�Wَ[%w��	�j����\���⏐U���̟���(�9�f5���27�ܤ�7����]�%�]Y`�M� ��]�;:�oҘ��Z=u蛟�tA%�UH�MA���U��Se�]8?i���a�s9o��ajr��OO��ax�K�wѪKU~L��[l�_��$����N��G�f*� 5IF�h�����1�����uf}��4]���tѕQ�33J���KG3$���؝<\C4b��Vgk����-���=I���o��S������N������dX��8]L�nխl�P����z,?�8�5Z�����WK��)`�y���f�⫦4���⸙�D�f�5�'YBz�3���"�3S�"��U3�@�ܸ/����>w
;��Ā?��{x�F�[��%S3���5��y�zFą�8�#�4��OW��@<�I�4p�&�k��S|_=	hs��fN�Ĕ��A��-+�gk��(��<�VWTW�βz���3Xa�e�tLůg>�R���̿b�ڪ�0�+��%�mU�f�S������
z�:�qZoA����z	:�T�*1¹�ƿHN�}�g��2 ���F��⁸��ր;g��^�4�A}�Ӛ�|}t�J��\�I��i=m"P�~�����b�\����_�,�Z��B
eFg6~�AmM-�����n�3b|˛��VW��ސ�4|�����7�����fG�����!�tj>d�UQJ��k#;��s%��ő���<"�|�D�����D~l���I�1���i
E�$���eY���E9�Ӹ'V��f�TjMzG�"u_?M��9Ih&`q��6q½�*|��� Q^>�5�h�3�J��L���g�5e�axh��Y�W�������V�X�G-ok�1z�B	'��rZQX�R��_I�%"W�w5Ց��(��W{���;�z��^�`�vT��}�p!������+"݅8؋vy	������~�zο��3��=��p1@���0P�_C0D�ಠ�X����;�?�ı��ۡ�!eԍ=C.�>�U�"���@�=�ar]�u�¢�ǦE��_�Ū� �e���z��=d�>w�W�� c��T��j�n��c;'�o�!�:yO�X���D6b���������J�]%�۬Oґd���}Pй�Of(�v�#t�)�����I�j���;gT�Ν��re���ѡo�~�'���n��v� �Y�e�Z�Q�@�"B J�$ғQ���-ƾ⯳ճ��*������b�4"M�A��G�bP�{K��������x�=��݁6��j�~N�Q��"�u�G������I�̷���^1�-��R�o��)	9�@KF��o�<�"��}Ͼ���k~ϛ�Ɋ�fv&���c�����t�̀uL�Z�(u�>'�mP�����N��fE'Zg�ӷU�/fuZ�Yj��w����� ;�5�71z�?=ϵUsm���Q=Tgy/Bz6�}��h��t�� �zEn�����������'�3�4���o-�3��W��_�M�)���(�3?n�;�@c.�m���b�����N���D$�mq��ȧ��bʱ��v���RN�`�f	2�f�''��[�ε&�G�n!���O+>��7�ƔFJ��T����0�
��X^D����ɓq��#'�*����O��Ҷ��p���\����dⁿ�i[L��Ӷ�Ò�(Dd��$�y,餫q����Z��#DO+4�|�s�o"C�^�b�DC����H3t6U�e�{�,���4���������S�|���O�����6Cv�Y(�>XDt�9����H�����m譃E��
�`��׎ ���Ym�S� Ȩ���x��h3�J�"�#�_�)�X�{���o� 1��~3�:����K�$��z�U
pGl��F\H9�[�����1�y��tHô�8���览����tnn��\''�7���H�]F>�m_���87����
2mu���UE[�����a����ځԨs\]���CF�ߘ��E%��](�x4���!�n�\YW��;Q��j��l�h�A���}�y��N�K��<��a&�'�c.�$A[��)��CLN~�b�f�*<�ڍ��m�$s?qh���1	$`;���ڔ�Z�B׍/	!ʠ˧} [%�h$] ��ĳ�<�sC`�\����-��
�K^7vX>�;��dX�^��U�M�f�zn�o�F(LYx2����f1KkY�F��W�����.�A�[2r�n�����\�8+?g�6�H[�RCRgh�u��{(�bg�`KE��������gRǫ���Gp�(���zyHz���V���M56��zu2OٽNqT/b�z5����a��8�>���^?K���ŵ�ϯ+3IH��Oy��]!�A��lB3e�h_�(� ��-�|�����Z�(�d���9����1�&ɏ�>w{���{I6K�Z	��+�f����sp߭8�	c����@`V+:FK�&C�mͬ�+k���.`be|���4-`V�@�ɬCd�XՕ8J�E�>�I~�<�F�3`���nR R��լ0��f��v�x�:Ѧ;�V甧+�'}'���U� /���8l��g��%�ٙ�~<_�+љ;i�Y�,�8u��/P���j��߲�e~Z:�X�^ ���ƪ���z��C��5�W� Y-r��w���%��:����ŧE����B�kP����O�����x�g7�2�
}vj��-=j�b
�w�{��J��,���
�VT_��GP�n6�l�R2�gi�L)~�r�!�Nx��B�v�S��b��H���"�gd��̋�"NYށ�pX^4�жo&��R�Gz��L���3��;V$%��֪�)y�������O���KK���I�ǅQ��z��q���1�8���4.�Z=dM�=i��N5 �?�&{�� Oʴ�N���6���x���7�tQ�0��9i`�C�H�km�ʮ���e�\��_��r���?�H���bt��J���7J��q��gC��x��}���S`F�m6���[���E�dix�:6>�6�ǻ�% �k3�iˑ�rC�<g��ӊ��yǨ�9;��"H\�V���y����;��dg�ٗtC���x}r/(D�Sh�����S�G�%<�nR�_F4��Ԙ�L��_���͟�$ �۪��r��ų����D�Zv"X�'.z����}���uz�J�_�~a\��0���z{����V��,=+�Ħ6�q/d�d?lm���x�NA��\��[��~
�T	E�(��\�Q�s��!'����RL��m�)yg�K�����,O�O�3Pr9��ߓ�AY􇔤f~5c�p32�ų���8��C�e�y�ޫ�#)3蕜��˂�r�p��t��?���"��|h��|�!�Ev�PrYCL���������q��7�p~b����	v�w
!�de��0_ì	�9��gL��bo�-Weƭ��
EN4�y�����W�de�-?Z�g�3�2T��j�����iS9�����x�h�=��_���n=t��e��=��AVM�e�ަ�����J5�p����L������͝�C�N�1<��th�2���g"w諯��"���f\��N.����Bыޘ<Ε��~5m|4�ù��u��t͈vډ5�x�fB1>bKө׫٘X�|6ו�?�\lV~�v��`�����{3����H1������_{ǃ�m���sj%[a��p
�e���n�W�36
<ֿs�Sx��Z;{�#�1��^���#��Pf �6s��u�;��i�lZ���o��{�j��~����,"�=���f�f��鳏��Ma�/����e��ƅ��o���P���V�f�ı�π�4[��D۔q�-xf^c$��6��M��l��FMV�Ը�|kF`��=��z+��C�k�KVN8�Y��)����A�zA(�9��Ox��|�5��L;U��`�5���o�E^�©+�=4g�NWLU�tW��K��/ݵ�32*���-y�9� �C�� ����tUU�6�riEh��R������x�8u���;r\1��~��x�W��t�_e��cFJ�y+
�	�)��4I�#f�9�������?0�����X&XRf�_;�W��T޸m��
rmb�CcE������wJ�������q	_��������[�~����$U�� �-j���*C����s�5�#>��UԸ베��q���S���{���^�h��nm�� �㰌~ҽHn���Xn���-Ӭ�z���,%	��\�h�y~�Eb'�'�-��F���d6r�f5��ż&���DV��Y�Vf_9ۃ��QZ�`GRo�������:I�����Q��WI�>)�O��i���+;i�;������M�G$��A�NR1�>��5�+? <q���@��w�a{����kj�_ۧon��&��Z� W|=����<�2�b�%g����b�K�b��ϗ��n-[o�A�L��/��5���t����^�B���;{u|��"�/�]��^<ߔ�5�;����ZS�[�����J��f�?��Da��"�隍XXULp50[���]��{��y�n�^���\�t�|�5����(P��ft�I�.t��p����	;��ujP=Ë1���$���Z{,�C����b=>���f��QYA:<����G�;�'�1q�����D�M��ך,7L�8��y��?j���$�!��T����BW�n۠���	C�N{}��𝭟�uQ�n&�J�ipF|wu�N��}<��fC��; Fs�=ʤI?����u-����>Lnk��>��~������Q���+Ӱ�wlA+x�Ў������3T�Z}�r�Y��Y�0��&�rS%�.�Y2��x5��G~ekOr��������j�xe�< *�O���rW�rЎ���;��D���V��V���6誓J�d`��$#�x5�g�XM�l��ٓ���n0�d.�S����V��/�.}Ÿ׊>Ύ�z�_~���O�����C�ֵXV���x[V��))oc`�%a^A�w3`�O��+X&��}+�x��Zzt6E��fT@I)���7�O&U"��j�[�lr:]�X����zm{�&���t�Q�l/����<�N��y��ͯl_yf;e=1���$�,�3��ü�ݿ�FD�
��a��Y5�����d�ǡ@�����us������i�ʙ�2dYCt�e�Ͽuno�n��KS!��)�5ÌH����h^!���%������^��$��>�c���E�[1�P�~��]�w<rx守i�	W��������\��.����y*r�mĳ�HQ�')|o0���m���$�Mʰ߃ܲ�D� �k�:Q4c�^�c�'=(���R\q1C*K7c�8�FP|{��L��~�=�b�t����,�o���c�k�\�YO���8�:/�_�R��P8uj3��~�F�z���Ǳ�]��� ΫGa��+Qn�7a����2��*.���~���7������l<��^��PͲ��'��O����t'�{��3H�ZA�a#����ih�L:Ej�q��fF��x��-n���>����Hr�1��6��u��t�PJgM�R+��l�bK�J\�Jf���1�o��rtT$8-\��=�����6��d���/\�%�+TH����r�yIUT2������p~|gqך3KW�@���i��?�8���Т��/��'������7(��t����+�6{r_>/���W}�h;�/����U,Qܘ�k7�����2&�F���	��#��3)s��qh��6���e:���t��0�w�Y�t��ڀ��Gm�K۠��ɭr��t��Ȇ�����
���J\������S���ߍT�n���,�:Z�\�x�d�UQ�M�d<R�e��0���i�8_	7���#�_�gl���vL�e��;p=I8����A:B�Dųf]�|&jD`z]��H�0-��OJ�0��~�!T�z+.=��y奉Z��g������>Xk�M
7I3��ICX�ZNWF����!��_��ت����� Y���2J7�eˀ45@N�n���2��>4[�B��O���i��پJ�b�2��M]1�t���6l,����-҇��s�Rd�h'�k'���Z;�$�ȏ�����걍���+������/����_8�{�\�D���s�t,uU�=��x	��*��Y��3v׬/���5�������W6���<�[,?i6�9�k?�?���V.#����؆��0��K�[�:�QP�=��ƞ�tO�RSy�ӄ`b�J��L���tn�K�noN�B2�Wr�Y���	6*J�ם�p��-�o�����m'�h-�{��Y7��9b$���#��|i.|}3�u~�!Y=>�W���|��6-$�ޖU	���.+Ÿ{q@������QԵ"���,,��ũ�aNwW��EX�!1��P$4z�#�7!�b�`��@��KWHۥ�`~���?yD ѕ�A/m��寙A���]�O��	��^�v��F�Ya�x����u8a$�1j��\�l�v�6�ΰ
b,�4ˊ�0�
70�5{��s���َ4~2��6�^��z$�`��%�ۀ����	��ݙmr����,�Q�j�Z��K;˗0y�0�4�:���u���@>�l��.�P�O��/��p[��/�:��'�0pO�j����B[9Ƿ�G*�5g���i\i4d��Dl` M�}кd(=�c�9`,[#K��U� }p!j�nu���׽���~��sk�0�����(�~R] -�)���@�[=�o�J�_Q��L1�-cf�B�8MhY�7'�GE8�D��V�-�@�H�WDF�A�Sb �)BkPμ�����l�!�։(D0�ђ�"��حh��oV������K�Q�Jc��p_� ֢	a�����ojV�q^Qeu�<u�"�~&0�g�-R��27�w��0)��#�k��M���濾JK�ҟ��e3'I�V��T��n1���2�yO~��W����C��ݸ!��f��$l7;��6�Lڣ{q/u��^?�� l-��T��i�r���k)SM%A�-�y	ct���M,�����J8)8�����[���vZ����j�!5�x���-���M���v��thCR�b�\�p!���4�z2)[�{�N��j�)O������z\��5��6���H��̎���H��֥Dߓ�jZ���H}�:��W����sk�.e�d�\�~����g�xi��/�Ľ���.�����1��*��(�XAE��tZ�i����)Y�v�6���wm�hFRǈ��q�U&���,� B�H���b������y�q�<\Y����a��YjGL�D�� 7��N�*$�����;�����bUs����V�A��;l����r�@��쳔�S�G܏+5�V�NZ�Oj��QpL�rP	��*5�~��Hx���v������;��z�����Y����KMX��Rub�.)����q�ty�$��e�'�Ç[
�|,��'/1�;3�Ι�^￥�cV�!yQ7=|���NH������yq��E*s�#ɇ���ۼ)��Mǯs���雑���/���>l�g�J�ե+7g�:q�:��)m���f�0n�'|zb���O����Jq�ʺ_��>��b*KX���>d�Z3j� 2
���
�s&n|�	��z����r��=���+TD��y�\������z�����:C������ª@jfFft�N'����;��xg8�Ҫi�;[3���LI�¯�Yi��؃tY�D�&.���\]��si[���\��Ii��<�XJ.�r6�i�Ο<�fU�S�F|�{U�ÿ�]�blĵ����s�j�!f������d�.:��mVo>{X����;�dW!�Č2���Ro��xM�ا{U.-�l�Y�AnV���+�f /玽��lÎ���PiӰ,,~�5�Պ�%� ���+�s�������]sK��W�WH��W�^D�I1h,��S���qAc��P�i�o��g����� ��̗�n��ʩ̷�qM�vl�ʜ����������X���|`�]�ZP��pg��=Z��=�$(>��l�7���Q��>��m�*Ġ�d5Y�/���?�b��\�����-z���YW��O9F��4Pj��1IҾF�2)�W�����)t�k�yaamR�|�
�(�G�m��I�7R�ٯI��3-���2�AA)�V�Vn�Gw��8]r�_�R�h�fkUK�x��Uutji�+�Ĺ��Mlv/n��|'�4>�2k���}V&&j��%s�u՝���،4��>�uzXKF${��]~`��@�4MJ��@�����Qt�oro��9��r��C����$��^H,�i.���>o�
3�T�	}DZQ�n^#N.C.ݔ�$�*Q��Kb���	h!䟚�O����'.�bN#7���#��eG�)
�g��V��tD+*���?��������O��x\��M���~\p`p˥�0� ]�:��'��J������t����e��ݯVK�"�	�^u�j���>o�`�镯!~#��ȳ9�"Of���ڟ�E��˖�1��B��4�҄9�`=7�U��.�R��v�s�f&a��z>0��-U�z0�2u�n)W�*M6ȕJ��Le7�5�����{>w�S�@�'/lƸ��c�	J�7·�v�?�U{����٫t���x��Az��2jS��ff��|�E��L3�c�d�=n�ы��
�z&e
������ɫ�6��.���c��W�A� ����
tF<(�jy�
BN�ϐ�4����OY ��I���N|e���F��H
?ޔi}j&����F�bM�����F��bΛ��d�>����b�k����eڴқ�>L-�nUg0��������[�2�T���t�>����+#��>�W�i�� vq
 ��Y�Y����<���倄bӲ�.�����궊��~_~�������6���2�������i�XK�[7�-�/_n��o {c��h����
��p:Y'0d!?��ǉ�^�jG���/i���ɑ�R"�K�1��~��*�_|��w�OjQa�P���fO�Iϙ��:c�5p��/⾽yq?L.?y:WL�%��V��Ì�(U�;I���" ��|�/���E
	k�Bt!����G��Pfs���"]��?�ٛK���eh���t�@��^͟hM3�Z�Qm�%�ӄ�P j��e�\%�v��у�0҃��^��)[�\D�0���H�WsO�(O�9���o(8*8侄�]��L(��=��#qD�`f�5�w
��(���!�g�o�I��	���'C�n��as���ҳL�g�%�p�A��-���:�D��V��:p=n�/���\WH���ڥ.6-nA~k~���K��~���PJ��)J�=j���O��Z�:�٠5�}��t�����~�(��KXcUplWQ�Z���?꓀��՚ܑ��� ] V�����|L��J~I�ѥ袤�^�E�
��Q/�����W���>�>W�~պ�ŬE��c2W��?�œ����vԻx���*����yZ+��z>��t����4~�o�X-h����7b�����^�VՒȝ:P���C��0w�sp�Q��]����G�*���p�ӏA���CU��E��S,l��%cuG�T��=|��u���5�4���g��'s�[��=W'�E�4f�'���7l���8�W��_3�,�Q1��6hϫ�d��&�� fҷQts���H���'����)8���7q��Z:51��^iN�_��4n��A!鴒}��6c��ll�S�����i\�'�/��DJ��P����F��o�ZM�µ+�9ga���T�f�Ş.Z�%��-F�T,��������F2��q��!x�[��-�$��湤���5�w���61�se�D<^r�߰<��B��u5��}��	KC�N�$2�<^�F��X�=�dbBE���^^�:`5Q�W:��C�������<��> ��;�>^�H�}Z�!��r�-^<=��剈+a+�o�'��Q(�V��������=3�+�ëi���;FHO)<c
.a�0�o�@�I|9�%�Z:g��x�笂f��.��ʝE}���&�ԃl�%m��a<�q��Q�ai%�#��i�C{��u"�u峿�R�R�����aMl[�Q��X! 5�HQ����JB��RUD:����D��J�I'�t�(U�.A)RE�$!��P�s�i��w�w���?�	ɞ={���[����kϭ��馤�m�pHh�K�`VC��yz�|�(D�c�@.�[N%�0g"������q*-`؜�$ot'2�_IҺ���;�gM�沁�Xuel���o^�ۜ`u�@��jUưS�k��A�����G%O_�FR����iߜa��g��a2�U�CDL5��n��l��u^���gĊ�E P`%�YSRwbٺ[�@Y<*���/x���ʧ��=����S6k�=>�y�cR�?�O�a#��vP5!������+�-�����0�����ϟq�R%&ꂜ�A�w�(W����Dת����*Pݻb��N��S�'�l֪�>-*���o=H�8��Ɔ�S\.J�U_�w�n�����b�\]5ˇ���N�M[��.�e�L�-n
YҮ�w���ic�z�:���^���s�>L�1��q���R��;��]y{_��U�g,v������OV�^��E���2�˶�
)8�'	I0���5�L���"g������6��4����(�!�!R�<ف8�	-Rh�_�YC�D�	��~�_q匢˞$K���H�S_?U&�N3�wW��_:xe�uzA��>}O����I���|��؏Ͽ���{:��$ibqi��؟�--�GF���&�9�0u��r�1���d?'V���?�.�)w�>�-O<�H�n�t'�|�����_>�y�r�ِ��1u���� º�<�Nrb��B����W���IG)I�t���/�Ą��z��ten��˱�1�+^�p������Ѣ[(_y�����).��O����k���I;=L�l^l/h0�D���BZ�x��[�d�lQ/�Zq�k[���������Ď�U�6	�=��m]=o��jI���~������S�~R�z�x�'ћ�A-I@���u�T_kP=�W�~� s8m[[�A�q���R�5$��� ������v/q)��=|�=|��<�1��Z��C�>"�Ֆ՘bA�����N��A�z�C_�Dl�ǿ	f��=��f%����.��Q9�"�{��p7�_�)�?�����k%���&�3�0�΁|�=:�
�GM8��Z�h�Є�Oь'F�
�dn7��g9$�����t�#��G��g�ʿJŬ0�h'q��ɤ⎂l��!J��س)+�ō� ���s�N�Q�`6:�B���H �͖|�g7�� N�Y�@{�YQ��yVt>���<dQ�2����]�K��<�+I���{�{�8�6��y8�Y�ԝ�l�IU�}߷ͷF��dWw�c�59���<K��a\��H�[9�V�xr|Y�S���L3�JQ~��z�T���V�.�'06z�:0M�~�&L�p�)��(�����w�4u�&�~�ײ����P��;J�BǷ�H;�`L���>�� ��Vt�V��X�w������c6%ίC2"r�"h$p��ha�s��/�w6��Z�"�Rݶ���,T��aoq���iM�o��,�N&���="Q0w��p��$j��Ӱ����E�=�!�]��O����'�8�҅��?�O���F���"h>a�|�u$���XS��=��{������-jړ+;�
�����K���1ﻃ�H�� �7���;�4�y�c]�x޸�f ��/�a��Z���r�v��]��p��K�xJ����G �!m���Ц�c�HoR�#���Gە��Cwqxf,��0~�Ts�6eO�⾇῅��:���O��Ph��J_V�ϝ�ne<O����F�~m��f�؝�Fh�4�4��R.�TS
�3S�w�e����}l�*�5W�0�]M�X�,�%������P=��ĲnJuH#���),�G��/�@�E�|z��]|������� ���YƤ=�qy�����Q�A?��I�~���V�7n���D
5��j�5�	ͥ~ų~�� 6�N�rx���g� 9GC��L�3�ְ�Kme��k+/��&�0�Q=�� �C��y���ӻOe�f��j���ؚ��۬��C=���^ut)n���lHGc���ϝ� }Hk��oFZ:��L`쭁-	�? �����_iI�=~%ϛ�)A���;A����%��e.�;)���s+�[�8�;�,K8����F�U)V1K}� �U|�2% �+v��(ArUb&w~d�^�!��Q���8��Ŗ�J��0�拨.���z�e-
�IN 5u��]g�@��]Y=i#�|�����L�kE�5)[=�cL��ƺ}Z���l�����[ ��L��|�A,�o������"��w>��v�BJkg�	�j�T%~9)�R�$r��(���z˥Xʨ�m��͆�}�C#ǳ���)}V� �2J����wi"l�����À�u�AR�߇��/S�@�t8��m�Tj�j����Od%��
(��r�J���Ц�Of&�z�����@��V,�#�Ag�z����`�8��&�!,�*���E"�h�H�5���{~M��P�|9�R��6�:UL�-�ΞzD�i�j4a�:&�J��J�C��
�<��s���������%�H�3��ri�]���m����$�{DSFN��y�/�:j����{4�։�"YiC��k^��p�xU ���w����a��ǀ�G\6�1�̮6�fL���zZ���g\M�vM�o<6�(�`�b�<&x����0��y(�6�K��Y��l�JD���9R�-t�eˬ�ˌ:H�v�3���=�����ٶ:��u��i�on�u�i9ڗl�4�|Nzv�)T�q��Vz����*��`(�vϽw�𤿵,��0m$s)��i�:�E�
����E���]�}�k�����j��5~9g��န���g��h?}�=v+��e�˳�2E�f5���>����!o�d�z�E�e�Ǻ�a��Y��Ӝ���o�{A������zx ���(],���$�|LSŊ�X���-�Я�௾�ϧe,�>ǔv��%�sk�@�{{�g�W>E7�*��9�{�R*����g���えw;���^g��pѵ-ȷDj�e��YՔd��sr�����-r�[���������
��2὘HcYT}��{���dV�O��t�T�*�j;�{}!:�K���]�]�A��g����t�8���I�6��?K�CK�����P�a�����O~W�]s��O1�:gXL/��寈 Ɂ��Y����Qg1�"�U���t�Z6�kz�mba�o����,iv��ê�"V�Nrf'��� ��R8`g��n��i<_��5Q{�9��X���	b���m��� ̤�� �ւTA�mP�@�-��8�6OpM�0��7�]e�����ei���@���|Br���㱉��������2	\͑$<b�t'�I�n�H+Y�K܋jfGKn�k�w�#�?�~�IO��R|���,cK�ޙ�6��<�#�iP���(��+Ǟ@Y~a�xJbo���oh2P2�ެ����\��w�������[�>N�0�� �ŏ�\� ��b*��t����01Χ*��j���c�>��P��f] Փh1Z����<�׳x�շ����؞M%���\E�f��w�����}��@��%1�A�5Ӱ��k�7O��:a���gٝ�b؟ڎ?E$�J��$�f��J]�"P�� à3�L��N3�'2|f�m���J��Cp���	=��޹F�J8��VC;���r�e��Z�|�}E\.��F��B�g�+�T��A�W��ۜmDbl-$1�՚�:�&�)d�!%����&�,- �\�򩁟�,!��l1���&3�vC���( �1e@C���>��H����\<xv�ΣTG�dJ����I� =�L��V����n�@}~.~�'<�ޙ{=��Rg���&mgn�k������m�Woh�Qu��m��oN/�[�T����o�+pA�ߴ�8p=�S��i�4Tǵ��[�M����m����ₚ�zAO>�߷���?1W���4�5��M�ˁ�1*d��{ I�ǡ��D�vOJŲx>#A������M7�2WP\�Tw7�a�9.��h�*mPv�����Jw�D����㒏8�aN��:����IW�ʑ�>z-���E{�&�K������ק�8.�(�9%9wAiC���(+�j>1\�Љ�y8s5��6Əm@�_rKt��m����\ �����1�c�y}�j+	\h��0TI4i#(� ʍ��y���U�w��[�Y�H��7�:�څ�1�C��gy�<ևS��g�L�d<�3�;�-+�j��߷2�~�'m����{j�-T��N�eR��>�Z�}���D#�������Ы��5�P��f���,P�����9�W\ƆeNi�D�;ߤ�G��?���ܢ��p�?�;C��ע�L�PT�R��hu�l�c_g�sɡ#���<
�s/���1����𽑔,1��_˰}Ћ�� ��@}�6�V!�k�MY�Go#�f2��S��$<��������O�T�[�*\e4�l"}�'ǆ9g�|�'{����ky?����j�G�;xgL)xN�MU/�N�3�Au�N�ݭ<cj�zxl\.j��K�	�:����RF��j#�JZ��:�Ȃ������S�T�}m5��k���ax'�B?���#�^���N�2՟�	!�hEZ�K?��R����u��}u؝c�H���F��>m:��q#����=i�sa�žVyU4�9)c�w}:)�:���|сuc��u(.�E�� E�4>��-�i��&MƖse?c�)4v�A�}Æ}��J���Ѱ����F������jųj�C9o��!�WYN�J�G����Z<��e�ڃ��/�Z?+4��p�gi�h�^�Q�B_���^ms�����h�k�݃���հ A>E��ca�ʵ�6���\��ZZE?��E@�6���/�^�rE��y~��1	�ٺ}��6�����|c����Â���!';�Ύ*��?��bԪP�=��jL��Nf��N���	Y�����n��vһCr���mXy�D�6iK�ýW?�b\�/8��(�i� 4ۅs$G7U�ɚ"ǂπ������P	H@�|NHg�Ǯ`��~�fhk�u$fM�<mOyۈ)� �F]�C9����}X���D��wذ�ÁS��H���P�Yl������KC��f�B���0� g>��^&����]���t�,SZ\��B�4]	��'����>5#���Ĭ(�}E�T��a\z���,N<�H�9f�5^;�?�	NKCdQp0��<���6�.N�E�h@������?`�[�s�5�?��ȕ�~�若���fꐑ�����7g�iT���%�ŕ���I��IһzF]L��|�F�G�e�[	���6�SP��!�F�S�J*r���+I�oRJ�l�����r��6���h��ݽ5QA�~�Oٖ)�f]����8,��rbB�5^��{�{_f�j���tپ�����ˑ�
��l%���1�_��6^E�\�i<���D�n>����i��o���xHx�wFy�?��wb|�޷���(5"�I�n��_&���$\L�3h��
�ȉW~(~Ć�� C�Rφ5�?��k^|��+�6�t�*�4�Z�3>��Gݽ�!�ƺ���Pk���{�7ݚ �$�ii����A�;D�wr;����/䁯���'���%�i�AhN�?jL �ւ�W���\._�9�5�%j��d)�{Ѭ����$�1D*G�#��Ã��/\K���)�����KK� ��3�k\vB#�tL[�����|؞̎��{��[!J��[��K�����3��Z����/�����83�g�l�f^���f�
�ذuDqs��>ږ�=:4h_'��b���R��j(�D�KF0�8�@3��^�� �hl[��y��#��'`���ǣ��.'�lǆ�	����
{̃�aD��)��0KT�U��Ӻd�7�ڋ�ڋ�c+�^��GM�E�ŝ�l7��)lX�Z#�	�����dj�`RG��7)9esĽ����,��7|���iFA�̊���+�r���M���G�߀�;>�wg� �N�<�഻�����=�d���gb�M"a��.�P�;;�:_�P|�W���G��J58R��r��}��Zq��=�ip\�)߻�v��F��'s���"hv�e�(��!�I.�~m֮��fm*2j��q�ֵm���a=x�>��r��hj[�VoX��������^�Cw:�c�^U[�#�]���!�l({�Dm߷��>q��ϥ��B����!���BY�<+�a�ߣ��0����s>H�#~�2�[���d	�7�eӋ�m�S�<�|F
�C���q���_]�A\�ġ���p"�Sr3<t��:�'o%f�|���/� D=��X�N)�獏'�9'\c<���TkG	��󟐶}�����Mr��!��*�0R0��5�<��![���?�[�qP�ֳy͹ђ����z����.�Tf����6u�w1���h.�ܖ.�T�������t����k�ѷ��K���y��GstQ�~g���q�����[���v�k6�մ���B����+���O����-?��f��e2�j�!��3�-���%DtMbA�k\JC SnA��y�"eX���)8E� J{ٍK�
���Ro�7��H����������n�$�-~'�><9�^�_�[r[�k)�f;̔��&>86H�����+�/��K�����:z���5����k��q/����sowg��پ&���p��)e1�x�4ChH������]vB` k�=�l��v��ޚ������I�VB^���ϭ�Ѡ`�����i^� �1�̐.�ۂW�BohgO����0�Sz��K�ۅ[�I����q�U��oR��O��\�2�u���>���<t��/��a�������j�Xf���L�������AAc"�9^D�-�7�w�o�2�C�~��^jʗ��/��w+Cf[C	.�-������˔#m��5]
�k͞P��ʫfy�WR<�n`��R�%���1��|��_�^Y�L"3��b����,p$ �j@e��}�f?��|'f\�8����0��ʨ����D�W���9,\�h�E�iD���t��QXu��k#i/a����a8`%�t<{�_��I�v��;��O=�Z �N�-(�f=����ԥx���C���F��Q#�u�=��}?�aXG"�q��0�v�eH�y����<v��g�2\˶�
%s���r�8�Z��6�8̎��5�6��TQwh������b4�*��i7�l����o:�j͗lA=3=`��u}W��]�p)m�����i	���\g�i�Ú����Vս�syd�0%_~N�u���Vq:�s^Jב�-F�߷5����tP�v�@i|�J��AJk�����|�,��0fU���\������/l���E������V���.��dX��{d�mӄ_2a���v��Q��E^<oh:�hj8ܧ����!RM<�xw}|�E�▱��k�._��N$�2������_+�
��v���k���b-���e��\gB�v}�M��Z\P�ƶ,sI�G���H/�}N�l���^gS�ǹ�S���$ګ��+���=3G��??�����V�<uV��77slx����辠�f��܊�W��!���Ǟn�/	��������X�ȃ���WX�Ň ,��U,��E+F����	�͊�3��6��g�m�f���|�sx�o�s�7�L����y������}����#��̇~d�2�'r����P__<��)�:^}+���E%��0��\��"8�MǼBp�W��T=-]��K�f��7�Cp�Uᆁ����C��M�5(Ne�l�
�Ճ�Ğ6ć`���Ү�����|�s$�
�	[����"RG�3��ԓ}�h��="�KX ��'U9�B$@Ɇu�c׋�e�bH$��1�m?:���1���0�"�x��L7��߂��zfD��Y��`���Ө�=��;�꬞��2'�c�7��q)�e��f����uV�p�_T-�����Ə#1G�W���ao�2��pӓlX���S��ԫ
4}�	�w8V��$	[��;�8]�]o�v�#�f�Uv{����d�?Hڎ�,�����$f��y��J_��}5��G�O������x��짱޼�$�"�k+@ ��໹�\�Ϊ@��l�jP�\�/��u�L:P3n��H0�P}x��q��Ah5�C-���̚��u���Ӄ���:����q]��]w�9Y�G�Ê *���K���E���+o���a4��q�Û�����Z �)-���w"@�w�x;y��W�e�E9�"ir�/�ǃ�]�h?������b��Ҧf�
E,��ֱRJ����$��
�m=	�S�S�.,��ix�'�;Vg���T8o{R�<�$PI��\3蓔��oi�ua���_��ĝ}v���&S@T�m�H�UBK$��y8hyyA���m��"�ڥ�d�!e'Xri��+JLc��N��N?;�r�3�O�6�j�%��3T��j����}ņ��ʌF嫆��V��������Se�X������N��h�Z`�������#�~7���]X���`�M�d�h��r��a���-)@��?��c�+q�A��g�9]tej�g�>xhx��Ne*�!Kc�a�f�� � �ku�k7�n�M�G��i>B>�7N�1�� Arǌ,�q]Q�܉/EL��Oc�������Œ)Q�	�돡��W#��0���`$�t�C��?�O�J<<��������:���Ӂ�ڋ@ �l��4U7-t�ci�a���������&��͗���0�ډ��X�����+��j	
��Z祊B1���܍�$�Jt;��/lX�F����X��mU�U�ת�Ϛ;�#;.�P�(�}�T��!pt7X��^τ�I�F|�vέ\.Byq-�:
�'�lQ�Q�����@��b&1]@�Xi@�k�唲̀���.Rz�l�0��6?dn6��6%0"���[%z$Ur'��L��"��wXB:�6w�$;��� �d��{�"�S����/�.1WJ|�w|A��/,r������XON��X�ĸk�
>��f�]q�w�&Ϩ�7m�[��)  ��\�<�v�]
�b��jJ��4Mv��Fb	_��;�ҹ������|܏�W�u��4Y��6� R�tm��Jr,��5�
��l7@ڋ��%�11db�C�,-wr���px_��w�Y���/���/u�8p�a��{uh�,AY�#�O�����'�q�LT~֓�:�tv��c��ո%�E���ܶk���~ђ�ߛ�6�؂��\ƕ�V�T��A�������gR�Q�M���;��\�����ڇ r��H"�8m��N�Ȳ�bt��֒3jt�O����K�t4���C&��n-IB����3��:�ʰS�6,57�WA���ZB�`�pJ1�T���+"�"�5��J��Bl�AR:��2� ��ӣf��RepP:��f���?��a��S���_��Rb�/�}����;��螷
�	��'�����{��A���R�z����YG�'ξ�d*ϡ��c������^ိ4�x}v;��P�wH��}# �~�X_��ʱa�{Q�1F,.�\�vxy���yj/�b��1�ʆ)�яU��\�bhfx��-�D%���.���d��,�{ӑu�3 i�b�rJ=�W�c��-Mzn��s��'�>J��EL5�
�eFO$$�Oԟ�������Y��:��W�b6(�<�V!i��Lj�Yʸls)�Q�[#�^�؅��T6ΌH�$���!{�A��L�����o�4��ٿ��� ����w�3��oy����O���0)u��\�Q�БgSȘ��czomK�>P���)��ճ��g�����U�5o��m�A��[�:~?�B,����鱉f,Q؛���v���u^��.��d�P'��LS�ib�q{>�}zSsv���+�6�D�����"�u��|F��������@'�̻�B�Ѓg`�攴��tV�8g�� �&�kn��5a�c�`�fbX6i�T�Qғħ�7��_�&��{����
�#�����U��
�1��B$��1:�pR��	���Ǚ(�[��JG��i��%7���>q��A�c�04��3�a�!s�?�f-��,��$���C3t(*X��V2a�`�,���񍱞y��BM�|`�8vD�o�?N�o��b�@���[�tu��6��D�+�z�"�z����~+Lb��7/@L�� #��t��p�_���� ��װ��]��T"���㜟H�z�fo]��=3M �#X��IM�]j�.��q�@'\z&�T&i�Ϗ�a{�/��O�}���ˬs�G\����i��Fk�Sɛ�@ri)��[@�ڧ.�e�<\�#��Ge��5�#� p��7y+���H�7���p9Ne ��͍9��)�=��=��J�f�qsZ�׸�hP[p��/�Z���+桴�GW&��Ѕn���킾?����Y[�X�6"�6����65��� �(�ȯ�������!|�k�<tO�N���*��ʹ�Ѩ��<�Em�h/"P��mwfw�����'hq���+�u�A�'QB�*(n2��=���t�w�[zdb�L��ݗ����t�Wfy��6�P�<���1�9��_�_՟^==��=Q��T����s{6qӹ/QbC�X���T.�0�sFZ�mfȹ�_����8�o�wtӡ�v����{Z\	I���މ���0y�뮲��(���G�j���A���bQE�j
l6^���r.�%�Oֽ�qt�������0);;�l�!��X�����ͷ��PX�]
���"�����gP��şfUE��0�D�e�2~� �f����Ĺ��J6`��P�Q�<�q%{"�4�a%3�`�0l��W�������b�*R�6�� �ܥ�g�@����{�2��@h^�bk����9�laȲo�,{[h�g���;���́R}�!l l��/ac�IƝQM��	"+����\�|u��>+�68�+'kr
����8�_��2��U1��!�R}��䯙64t�,b�3��A��*Jc�92o�K�m��k׿0J]w~��bV��}@`����@9�&�˓��A�;��J{��͏Ė68�;^�?��l�	�jL��]T?TWt����4���Qர1�.�&���[�Y$�PTaN=���,KSD�U��T��LncB��T�'��1��0�uKK�M��&��ˉъ8�ㆣ���J4�7�82l[���A���<��3�����zh?���ސ����1Ȓ�m��!��Z�a� ��K{��f |���4�Q�OQDnG�g�D�B���)V�1�(%<��F�}#����������8�W��.j�5��8�g2�,�A�$~��I���C^�D�BG��݌[�FO�֜C�Q��-��&�3�����s��N�'w��h��)�o4R�[��_��^=�N%������?��b�w����yO�)��Glت	wz�rt��Jb�2���e����7l8��nL,v���)T1��Ӵ�x���sŽ���#G6�0�t��B&��ߚ�A}��9��|T[95�ݧ�sS������w���م�zl������E��)��O��U�]�B���r�SOCr�5��'�:b���Nm{&��Y�4����)!C�/�+�$�o�a�SB±a�fAA8�������V�
�5ԇ0���� x��ԍځԳ�WÃ��6K��<�g��w�ւ�*-�������4I��t���͸l/COib#����y����!���~k=kmH��F�~ω�c��I.-���Q��I2}:<w�
��z�dZFʗpܚd�?'v�1�렼��
[�"��f�O.2�*��8EB>��b��(̗$?K��w嶛ε�&F)\�'Ǎ.
�M�] �E6L�G���8�%����8>W6���ˆ��ˑF�g��1h��M:̓5�X3��f�����l~�	hf���k��,��%^G�G<����G"6���:ZR�뺵����6��(uOk�[5|�:ﶄ�B�i~6����>?�ž7�
@�c ��b 2��JD_�6KD��b���TO	��+<4& CS��_/-��>���!ؖIe�����b;��<�S��,�rC�������ߖ`���|U��'ݻ��Ĭi����|�@����Vf˰�5�J��;�~�5-�	��
U��܊�
#p�8LṒ[b��S+2������,G����f��|�43�.N��m�{1?�l�V>,�!k䪾�K;0w}��[l�_fEL��UK8�ʫ��~\u��x��؅w��ޤ�;&��6�Q���kD�Ol���4��Yڴ?��X���W�\��m`h������+$�k4e�άs)�~��p2|�%���w�~_^���~I��j�Q3����B�i���| e��ԏxnl��S[ݜt�O�Ӯ{"k�{r��}M�z�eGG��۟���P/.�s��P�(Ȝ��[���{�3q"+i��t�"��H#V-�k5��;K��Y�s��\��!H(T���
l�zN�i�S�$�|�"u�E�fVZ�A��~4��J�;r?�Df��r��\e��9��dbz��� lH�*�����`�����,��&I~���Υ�*[�����ް+��-{��w����G�#c#R�^�ċ}&�o"��'���H�Ӈ�g]�ˆu�zI\kbZ�a���ZM�'m��H�l"g]���ŨTA�������d7�������N�ǹ�\U���=e�үBrF��]J��M�K�Ⱦ,_w���g�
f+o9�X�8^yǛ���|/��!��m�A*��Fj�id"��=��T$�a��,��Vd��9��J��t⡀�h�֜�W���"�_�9�(O#	i�̘��Ĝ�֬��e�|����爋8���i�oyr����F�	���ؤV��w���w!��Q4�ٜ��X��,�����oc�����sڲ95�2��7�9����Q�5�f�>�^�0�怾������u�/4e�apV��-�K?�0-S�L� �Nv�ێE��}�����!n�Gغ��bF�.k����̶��ҍ�7� Ǟo�~ԟ�g�D�Es7o�ި/(IxwJ�HSD���hw��ұ�?�fS�HN�%�񽊸l�>���sX�;?�k�ZZF�e�JV�4�x��� �;�ְ�x�8�""����x�����"��s���׻X�i�&J�o'ua^̬�O�3$,���f ��C�4P� �W`��B��B��av�����Ec٣z��6L�PB�����m�a��7�ζK�uz��ܗ��<ˏf���)�H´g��Ð�ɸ�1A��D�˜�,<���Ko��~��^E!��*��hո�6��h9��h[C��b�P[eӫ����=V�0�xt�1p�gD�h)�>瑯��E��6����D�}bia�����D�w�y[�FX�e|óW��1|��>S�$���o��&���;�AZZGل�[K�J���S����tlH�%���_���<\	4�	���Z~�$|��Z
�kTUZx�.��Y��f�!�>'|P�&�������l�ޕax���2
����n�iS$N�fR`�4�/d�'7���Z��yB�qɢH�n���C��S)u',փԭz4tL��W�^�1�k���&e��O��v��ܽT;rJ��鐜��gK�&��D�DX�FtӶ�Pg���X���-���-�"s����BS[8��lg�v*����ď��`��p��������x9�N���nL��G��J ��&�E>�� � �5_��R�T�R^�'PO����Z�X�d�U���&�/���՞vcԕwˁ����g�޸w�4vCK�ڻoSuv��WM�_����Pg�s21��0W�'�����³���ذ��;�VxZx<�~F�g���&U�㧊ng�f�n4ɧ�����X�����F�HV�&9�d�E%L)lY���;��H�7���*`��}��UE��v$F�^�wm���s�MC3���C���ORٰs�����}�V�+��yi�q$Xu�Z�bu��Sn��ё+�s_O�+{ȣjr�k>s��5�IqX投����O%�m�0pv;{�N�}�<l)]�BDG�G�[��$�Ojf��6G~VA
��}��4�[�ȱ��5�T=R�[W�A|��n[S��=u��k�g�#h��S��/4?|e�G羐ZB#����.:!*1�X�.$4�A3r�V�if�H�?d��-��J�E�A���/�f���|��a%u����3�h����������������������V�c��&6,���z���;K���aE�#۷&�޷�aCbl]�_�.���Hm�$���ߕhΝk7��Q[h�ùR�KO%���!ɠ/��j���K��t��4M�B��+)������"fy�T��Vww��և�Q,�pz�Ӣs����y.7��Nr�Q�5�@� !�w݈R��@%�<�D��4!�VM��ʍ��uA�6F�J�I,z�YG����o�r?�p[�M��A��K�r�
�f��V�+Q�nΧ��<���D/l�m t[�HC@C�l�����R����/������'�O��B�؏�5/|��&\�G6���{�=����XH~��{e㙾��m�/4?x�fʴs�����{Cz��O����M=�v{F��ͥ��ǒG?��V���ݔ��88Y3B
�n�?PK   �N�X���8J	  �O     jsons/user_defined.json�Z�n���A}i=���tl�0�8���S���\62�PTr� �ޡ����I�@��z�iq�=�Yk�Y�����܍O�˅+�[����d�ŕ����?`�,�i�����_߷\���۹.?�X棛�K� A�7٬��1+g��J�?�*�]�E�-�����|�n��~�	~��l�&�,|#�"��R�)��@@t���e�}r�na�l^�3�_��L��h̝C���(����K�-�0�*M���p�<�/s_�O�����y������bF?�	�?�W��_� �3�̳�ː@~io�2�aJ�����U6W��['x�-�&[Ls�(���Ӫ\�I����7ܢ��qtԂ�b�9�����<��[�;¿=;�x����[=�7���5+���.��ܕU�YǛſXOt����y�=[����UX��2�6K�c��u~V��w��U�6[d�����r|� �A�b�|鵩��+��p�b��L��� YjR�	��B@�4@s�@�f=#T	�!�	q����ۭ(��t�?��E ��l��u��h�ѭ�BLK���bt�����LY���������� ��N=p�Q�U��S"�%�JvU�3
��������;��q�� �9��z��Ky��Ҧ�B ��_6�~�8����p�N����@��Y�����M�);|������M���n�m�F�����(8�����$
���#8���(��͢�2�-;b�(��b���"N�8Qc<}.��q�ve����9ڑ��a�Q�8C;���W�o/�!�4��R�O^]޾��h��?���˫8~�����	jR�?��&qy_)fo��M��Z<��7�����4.<��_�W��q��M�<��=n2����i�P�&yyOU��k,n�mG�N�+��ڎ��ƕ�p�#e�7/��-��HX����0��,��۳ě�&k�V�^���j��������M>��n����
�j��z>{ō��;uW�{n
�;�u���)��p�B|4����:�~�	�پ?���D�0�@�K�O� �B�{>��l�������zY͗U��Z��w(�!��R���������v��"�QG !ȇ13$�x��O�֘��	��]��tY]�a���Jp�!Qumq�=���Z�a��V*��,�DF��c[&��3ٖ���Q�Ne��5��.�q�6�B��l�+��z�>���kpj�/�Y5���'���e�J��e��:M�Oxd<�ʄn�:0t`��Ё�C5C�J����������Q����|����JS&���G���0<c�1z�J@39���eލ+ɕ�(�[1PXZ.���ͤ�g�A��J�(�8�@�JD�!H�9���e�ڏ�HX�j]�,�R1�}~'d��GL(&�j寵HD���@GB$�q��J� 
?������B�k|Bh����{�v����ě�	��������$tL"s�����i�ݳńu�o=�hڋ��GDu��˛��F�`��>�۩ɑ�<�a"Gd*�Q��S:'���+r��QF�e��ulU��[�ae.�B�B���G�Ʋ�kӕ��M�B�I�E)	�
�@� �E��W,�����b�*����dQH*��`ʓP��#/<��<�DœP��8ޭt�-���|�$ߤ�B��l6��^�N��K���lS��10�PJ���ء>�!܋�N�$�S��o*Y-�*!&������C��XS��x��C����#�⧐��}���;Dhy���m�xP&&&*PO2.�<���ϑw�!d����������dK@M�����2;�~o�������]3sZKk\�`yhFEh���X#�Wk��ј��]s���4� �2P�BL	`�q�S�|���=?욽R�{��,���;�:��aK.��Ě�MO�A2	Ox�J���W�
�Q�k��	S,�[��P�ʰ��1�F?ҹ"��Ob9&�b���>rH���?;'G�ȷب3�����S�d{@���"P�͞
�_�i��&J��@i'�� �5%�c�6}J� AΉ���N9 \j�7��}��zŏf�̪ok��	�e?![ˣrV���s�W[,0��|U��٬�ہ��Wv��ݻ��Tg���O�~��϶z���x����M�R؇N����,��jTܷw��b��6�c����
���g���ʤ�}��E^�f�q���O����Y�,�Pۮ�׶dmS�mmոP�B9�.�n'��T��^���<΃���a8���������<�q�lÞmس����>|�<�y������>|�<�y�����>���_PK
   �N�X�)��E  D                  cirkitFile.jsonPK
   �D�Xf�� w ߀ /             r  images/04914e81-76ea-41b3-8036-a4ddbf8d15ca.pngPK
   �n~X?�]��  z�  /             ߓ images/0769869c-6d33-46eb-8102-928d675c2604.pngPK
   �N�XWC��)�  � /             �# images/093f54e3-331f-4155-80d0-fca9fbcaa25c.pngPK
   |G�X�v��f �� /             +� images/153184b0-233d-45e0-a203-5756afb39f29.jpgPK
   �N�X����7  �  /             l_ images/2b66d102-ef9e-4dde-8ee7-817842500f7b.pngPK
   �N�Xo�>��q  �q  /             �p images/2cd737db-51bc-41eb-8762-f3273c40eae5.pngPK
   �D�X���(5  #5  /             � images/50d22222-f918-4c14-b9d3-6f9cf2edfac2.pngPK
   �N�X��_8
  3
  /             | images/57489f55-55cc-4ea4-8258-f1cf3d9c722d.pngPK
   �N�X�E��    /             # images/85bcb663-dfd0-4f8c-a6ae-bb35df534978.pngPK
   �N�XN�v4	� m� /             �6 images/91e5cd07-2a88-4b0d-9128-72e2f992e16c.pngPK
   �N�X�&�}[  y`  /             (�	 images/982accd3-ee7b-437c-8e9e-7ebd1fcbf7fd.pngPK
   �N�X��!O uq /             �J
 images/ca26ee1a-c8ec-49c9-93c2-f85ad300bf9b.pngPK
   �n~X����}  �}  /             O� images/e0206f85-8494-42b8-8b98-142c319be1e7.pngPK
   |G�XEm��O �� /             y images/f99a6fc2-4a50-4dfe-be0a-52d397e863dc.jpgPK
   �N�X���8J	  �O               �g jsons/user_defined.jsonPK      �  \q   